// ECE385.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ECE385 (
		input  wire        clk_clk,                //             clk.clk
		output wire        eth0_mdio_mdc,          //       eth0_mdio.mdc
		input  wire        eth0_mdio_mdio_in,      //                .mdio_in
		output wire        eth0_mdio_mdio_out,     //                .mdio_out
		output wire        eth0_mdio_mdio_oen,     //                .mdio_oen
		input  wire [4:0]  eth0_mdio_phy_addr,     //                .phy_addr
		output wire        eth1_mdio_mdc,          //       eth1_mdio.mdc
		input  wire        eth1_mdio_mdio_in,      //                .mdio_in
		output wire        eth1_mdio_mdio_out,     //                .mdio_out
		output wire        eth1_mdio_mdio_oen,     //                .mdio_oen
		input  wire [4:0]  eth1_mdio_phy_addr,     //                .phy_addr
		output wire        eth_pll_125_clk,        //     eth_pll_125.clk
		output wire        eth_pll_25_clk,         //      eth_pll_25.clk
		output wire        eth_pll_2_5_clk,        //     eth_pll_2_5.clk
		output wire [31:0] io_hex_export,          //          io_hex.export
		input  wire [3:0]  io_keys_export,         //         io_keys.export
		output wire [8:0]  io_led_green_export,    //    io_led_green.export
		output wire [17:0] io_led_red_export,      //      io_led_red.export
		input  wire [17:0] io_switches_export,     //     io_switches.export
		output wire [7:0]  keycode_export,         //         keycode.export
		output wire        nios2_pll_sdram_clk,    // nios2_pll_sdram.clk
		output wire [1:0]  otg_hpi_address_export, // otg_hpi_address.export
		output wire        otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,  //                .out_port
		output wire        otg_hpi_r_export,       //       otg_hpi_r.export
		output wire        otg_hpi_reset_export,   //   otg_hpi_reset.export
		output wire        otg_hpi_w_export,       //       otg_hpi_w.export
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire [12:0] sdram_addr,             //           sdram.addr
		output wire [1:0]  sdram_ba,               //                .ba
		output wire        sdram_cas_n,            //                .cas_n
		output wire        sdram_cke,              //                .cke
		output wire        sdram_cs_n,             //                .cs_n
		inout  wire [31:0] sdram_dq,               //                .dq
		output wire [3:0]  sdram_dqm,              //                .dqm
		output wire        sdram_ras_n,            //                .ras_n
		output wire        sdram_we_n              //                .we_n
	);

	wire         nios2_pll_c0_clk;                                                // nios2_pll:c0 -> [eth0_mdio:clk, eth1_mdio:clk, io_hex:clk, io_keys:clk, io_led_green:clk, io_led_red:clk, io_switches:clk, irq_mapper:clk, keycode:clk, mm_interconnect_0:nios2_pll_c0_clk, nios2_cpu:clk, nios2_jtag_uart:clk, nios2_onchip_mem:clk, nios2_sysid:clock, nios2_timer:clk, otg_hpi_address:clk, otg_hpi_cs:clk, otg_hpi_data:clk, otg_hpi_r:clk, otg_hpi_reset:clk, otg_hpi_w:clk, rst_controller:clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] nios2_cpu_data_master_readdata;                                  // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                               // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                               // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [27:0] nios2_cpu_data_master_address;                                   // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                                // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                      // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_write;                                     // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                 // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                           // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [27:0] nios2_cpu_instruction_master_address;                            // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                               // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_chipselect -> nios2_jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_readdata;    // nios2_jtag_uart:av_readdata -> mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_waitrequest; // nios2_jtag_uart:av_waitrequest -> mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_address -> nios2_jtag_uart:av_address
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_read -> nios2_jtag_uart:av_read_n
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_write -> nios2_jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_writedata -> nios2_jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_eth0_mdio_avalon_slave_readdata;               // eth0_mdio:avalon_slave_readdata -> mm_interconnect_0:eth0_mdio_avalon_slave_readdata
	wire         mm_interconnect_0_eth0_mdio_avalon_slave_waitrequest;            // eth0_mdio:avalon_slave_waitrequest -> mm_interconnect_0:eth0_mdio_avalon_slave_waitrequest
	wire   [4:0] mm_interconnect_0_eth0_mdio_avalon_slave_address;                // mm_interconnect_0:eth0_mdio_avalon_slave_address -> eth0_mdio:avalon_slave_address
	wire         mm_interconnect_0_eth0_mdio_avalon_slave_read;                   // mm_interconnect_0:eth0_mdio_avalon_slave_read -> eth0_mdio:avalon_slave_read
	wire         mm_interconnect_0_eth0_mdio_avalon_slave_write;                  // mm_interconnect_0:eth0_mdio_avalon_slave_write -> eth0_mdio:avalon_slave_write
	wire  [31:0] mm_interconnect_0_eth0_mdio_avalon_slave_writedata;              // mm_interconnect_0:eth0_mdio_avalon_slave_writedata -> eth0_mdio:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_eth1_mdio_avalon_slave_readdata;               // eth1_mdio:avalon_slave_readdata -> mm_interconnect_0:eth1_mdio_avalon_slave_readdata
	wire         mm_interconnect_0_eth1_mdio_avalon_slave_waitrequest;            // eth1_mdio:avalon_slave_waitrequest -> mm_interconnect_0:eth1_mdio_avalon_slave_waitrequest
	wire   [4:0] mm_interconnect_0_eth1_mdio_avalon_slave_address;                // mm_interconnect_0:eth1_mdio_avalon_slave_address -> eth1_mdio:avalon_slave_address
	wire         mm_interconnect_0_eth1_mdio_avalon_slave_read;                   // mm_interconnect_0:eth1_mdio_avalon_slave_read -> eth1_mdio:avalon_slave_read
	wire         mm_interconnect_0_eth1_mdio_avalon_slave_write;                  // mm_interconnect_0:eth1_mdio_avalon_slave_write -> eth1_mdio:avalon_slave_write
	wire  [31:0] mm_interconnect_0_eth1_mdio_avalon_slave_writedata;              // mm_interconnect_0:eth1_mdio_avalon_slave_writedata -> eth1_mdio:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_nios2_sysid_control_slave_readdata;            // nios2_sysid:readdata -> mm_interconnect_0:nios2_sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_nios2_sysid_control_slave_address;             // mm_interconnect_0:nios2_sysid_control_slave_address -> nios2_sysid:address
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;            // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;         // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;             // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;                // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;               // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_nios2_pll_pll_slave_readdata;                  // nios2_pll:readdata -> mm_interconnect_0:nios2_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_nios2_pll_pll_slave_address;                   // mm_interconnect_0:nios2_pll_pll_slave_address -> nios2_pll:address
	wire         mm_interconnect_0_nios2_pll_pll_slave_read;                      // mm_interconnect_0:nios2_pll_pll_slave_read -> nios2_pll:read
	wire         mm_interconnect_0_nios2_pll_pll_slave_write;                     // mm_interconnect_0:nios2_pll_pll_slave_write -> nios2_pll:write
	wire  [31:0] mm_interconnect_0_nios2_pll_pll_slave_writedata;                 // mm_interconnect_0:nios2_pll_pll_slave_writedata -> nios2_pll:writedata
	wire  [31:0] mm_interconnect_0_eth_pll_pll_slave_readdata;                    // eth_pll:readdata -> mm_interconnect_0:eth_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_eth_pll_pll_slave_address;                     // mm_interconnect_0:eth_pll_pll_slave_address -> eth_pll:address
	wire         mm_interconnect_0_eth_pll_pll_slave_read;                        // mm_interconnect_0:eth_pll_pll_slave_read -> eth_pll:read
	wire         mm_interconnect_0_eth_pll_pll_slave_write;                       // mm_interconnect_0:eth_pll_pll_slave_write -> eth_pll:write
	wire  [31:0] mm_interconnect_0_eth_pll_pll_slave_writedata;                   // mm_interconnect_0:eth_pll_pll_slave_writedata -> eth_pll:writedata
	wire         mm_interconnect_0_nios2_onchip_mem_s1_chipselect;                // mm_interconnect_0:nios2_onchip_mem_s1_chipselect -> nios2_onchip_mem:chipselect
	wire  [31:0] mm_interconnect_0_nios2_onchip_mem_s1_readdata;                  // nios2_onchip_mem:readdata -> mm_interconnect_0:nios2_onchip_mem_s1_readdata
	wire   [1:0] mm_interconnect_0_nios2_onchip_mem_s1_address;                   // mm_interconnect_0:nios2_onchip_mem_s1_address -> nios2_onchip_mem:address
	wire   [3:0] mm_interconnect_0_nios2_onchip_mem_s1_byteenable;                // mm_interconnect_0:nios2_onchip_mem_s1_byteenable -> nios2_onchip_mem:byteenable
	wire         mm_interconnect_0_nios2_onchip_mem_s1_write;                     // mm_interconnect_0:nios2_onchip_mem_s1_write -> nios2_onchip_mem:write
	wire  [31:0] mm_interconnect_0_nios2_onchip_mem_s1_writedata;                 // mm_interconnect_0:nios2_onchip_mem_s1_writedata -> nios2_onchip_mem:writedata
	wire         mm_interconnect_0_nios2_onchip_mem_s1_clken;                     // mm_interconnect_0:nios2_onchip_mem_s1_clken -> nios2_onchip_mem:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                           // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                             // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                          // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                              // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                 // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                           // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                        // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                            // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_keycode_s1_chipselect;                         // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                           // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                            // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                              // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                          // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;                 // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;                   // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                    // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                      // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;                  // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                    // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                      // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                       // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                         // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                     // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                       // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                         // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                          // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                            // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                        // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                       // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                         // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                          // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                            // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                        // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                      // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                        // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                         // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                           // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                       // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;                   // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;                     // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                      // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                        // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;                    // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire         mm_interconnect_0_io_led_red_s1_chipselect;                      // mm_interconnect_0:io_led_red_s1_chipselect -> io_led_red:chipselect
	wire  [31:0] mm_interconnect_0_io_led_red_s1_readdata;                        // io_led_red:readdata -> mm_interconnect_0:io_led_red_s1_readdata
	wire   [2:0] mm_interconnect_0_io_led_red_s1_address;                         // mm_interconnect_0:io_led_red_s1_address -> io_led_red:address
	wire         mm_interconnect_0_io_led_red_s1_write;                           // mm_interconnect_0:io_led_red_s1_write -> io_led_red:write_n
	wire  [31:0] mm_interconnect_0_io_led_red_s1_writedata;                       // mm_interconnect_0:io_led_red_s1_writedata -> io_led_red:writedata
	wire         mm_interconnect_0_nios2_timer_s1_chipselect;                     // mm_interconnect_0:nios2_timer_s1_chipselect -> nios2_timer:chipselect
	wire  [15:0] mm_interconnect_0_nios2_timer_s1_readdata;                       // nios2_timer:readdata -> mm_interconnect_0:nios2_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_nios2_timer_s1_address;                        // mm_interconnect_0:nios2_timer_s1_address -> nios2_timer:address
	wire         mm_interconnect_0_nios2_timer_s1_write;                          // mm_interconnect_0:nios2_timer_s1_write -> nios2_timer:write_n
	wire  [15:0] mm_interconnect_0_nios2_timer_s1_writedata;                      // mm_interconnect_0:nios2_timer_s1_writedata -> nios2_timer:writedata
	wire  [31:0] mm_interconnect_0_io_keys_s1_readdata;                           // io_keys:readdata -> mm_interconnect_0:io_keys_s1_readdata
	wire   [1:0] mm_interconnect_0_io_keys_s1_address;                            // mm_interconnect_0:io_keys_s1_address -> io_keys:address
	wire  [31:0] mm_interconnect_0_io_switches_s1_readdata;                       // io_switches:readdata -> mm_interconnect_0:io_switches_s1_readdata
	wire   [1:0] mm_interconnect_0_io_switches_s1_address;                        // mm_interconnect_0:io_switches_s1_address -> io_switches:address
	wire         mm_interconnect_0_io_led_green_s1_chipselect;                    // mm_interconnect_0:io_led_green_s1_chipselect -> io_led_green:chipselect
	wire  [31:0] mm_interconnect_0_io_led_green_s1_readdata;                      // io_led_green:readdata -> mm_interconnect_0:io_led_green_s1_readdata
	wire   [2:0] mm_interconnect_0_io_led_green_s1_address;                       // mm_interconnect_0:io_led_green_s1_address -> io_led_green:address
	wire         mm_interconnect_0_io_led_green_s1_write;                         // mm_interconnect_0:io_led_green_s1_write -> io_led_green:write_n
	wire  [31:0] mm_interconnect_0_io_led_green_s1_writedata;                     // mm_interconnect_0:io_led_green_s1_writedata -> io_led_green:writedata
	wire         mm_interconnect_0_io_hex_s1_chipselect;                          // mm_interconnect_0:io_hex_s1_chipselect -> io_hex:chipselect
	wire  [31:0] mm_interconnect_0_io_hex_s1_readdata;                            // io_hex:readdata -> mm_interconnect_0:io_hex_s1_readdata
	wire   [2:0] mm_interconnect_0_io_hex_s1_address;                             // mm_interconnect_0:io_hex_s1_address -> io_hex:address
	wire         mm_interconnect_0_io_hex_s1_write;                               // mm_interconnect_0:io_hex_s1_write -> io_hex:write_n
	wire  [31:0] mm_interconnect_0_io_hex_s1_writedata;                           // mm_interconnect_0:io_hex_s1_writedata -> io_hex:writedata
	wire         irq_mapper_receiver0_irq;                                        // nios2_jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                        // nios2_timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_cpu_irq_irq;                                               // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [eth0_mdio:reset, eth1_mdio:reset, io_hex:reset_n, io_keys:reset_n, io_led_green:reset_n, io_led_red:reset_n, io_switches:reset_n, keycode:reset_n, mm_interconnect_0:nios2_jtag_uart_reset_reset_bridge_in_reset_reset, nios2_jtag_uart:rst_n, nios2_onchip_mem:reset, nios2_sysid:reset_n, nios2_timer:reset_n, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                              // rst_controller:reset_req -> [nios2_onchip_mem:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [eth_pll:reset, mm_interconnect_0:nios2_pll_inclk_interface_reset_reset_bridge_in_reset_reset, nios2_pll:reset]
	wire         rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                          // rst_controller_002:reset_req -> [nios2_cpu:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_cpu_debug_reset_request_reset;                             // nios2_cpu:debug_reset_request -> rst_controller_002:reset_in1

	lantian_mdio #(
		.CLOCK_DIVIDER (40)
	) eth0_mdio (
		.avalon_slave_address     (mm_interconnect_0_eth0_mdio_avalon_slave_address),     // avalon_slave.address
		.avalon_slave_read        (mm_interconnect_0_eth0_mdio_avalon_slave_read),        //             .read
		.avalon_slave_write       (mm_interconnect_0_eth0_mdio_avalon_slave_write),       //             .write
		.avalon_slave_readdata    (mm_interconnect_0_eth0_mdio_avalon_slave_readdata),    //             .readdata
		.avalon_slave_writedata   (mm_interconnect_0_eth0_mdio_avalon_slave_writedata),   //             .writedata
		.avalon_slave_waitrequest (mm_interconnect_0_eth0_mdio_avalon_slave_waitrequest), //             .waitrequest
		.mdc                      (eth0_mdio_mdc),                                        //         mdio.mdc
		.mdio_in                  (eth0_mdio_mdio_in),                                    //             .mdio_in
		.mdio_out                 (eth0_mdio_mdio_out),                                   //             .mdio_out
		.mdio_oen                 (eth0_mdio_mdio_oen),                                   //             .mdio_oen
		.phy_addr                 (eth0_mdio_phy_addr),                                   //             .phy_addr
		.reset                    (rst_controller_reset_out_reset),                       //        reset.reset
		.clk                      (nios2_pll_c0_clk)                                      //          clk.clk
	);

	lantian_mdio #(
		.CLOCK_DIVIDER (40)
	) eth1_mdio (
		.avalon_slave_address     (mm_interconnect_0_eth1_mdio_avalon_slave_address),     // avalon_slave.address
		.avalon_slave_read        (mm_interconnect_0_eth1_mdio_avalon_slave_read),        //             .read
		.avalon_slave_write       (mm_interconnect_0_eth1_mdio_avalon_slave_write),       //             .write
		.avalon_slave_readdata    (mm_interconnect_0_eth1_mdio_avalon_slave_readdata),    //             .readdata
		.avalon_slave_writedata   (mm_interconnect_0_eth1_mdio_avalon_slave_writedata),   //             .writedata
		.avalon_slave_waitrequest (mm_interconnect_0_eth1_mdio_avalon_slave_waitrequest), //             .waitrequest
		.mdc                      (eth1_mdio_mdc),                                        //         mdio.mdc
		.mdio_in                  (eth1_mdio_mdio_in),                                    //             .mdio_in
		.mdio_out                 (eth1_mdio_mdio_out),                                   //             .mdio_out
		.mdio_oen                 (eth1_mdio_mdio_oen),                                   //             .mdio_oen
		.phy_addr                 (eth1_mdio_phy_addr),                                   //             .phy_addr
		.reset                    (rst_controller_reset_out_reset),                       //        reset.reset
		.clk                      (nios2_pll_c0_clk)                                      //          clk.clk
	);

	ECE385_eth_pll eth_pll (
		.clk                (clk_clk),                                       //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),            // inclk_interface_reset.reset
		.read               (mm_interconnect_0_eth_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_eth_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_eth_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_eth_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_eth_pll_pll_slave_writedata), //                      .writedata
		.inclk0             (clk_clk),                                       //                inclk0.clk
		.c0                 (eth_pll_125_clk),                               //                    c0.clk
		.c1                 (eth_pll_25_clk),                                //                    c1.clk
		.c2                 (eth_pll_2_5_clk),                               //                    c2.clk
		.c3                 (),                                              //                    c3.clk
		.scandone           (),                                              //           (terminated)
		.scandataout        (),                                              //           (terminated)
		.areset             (1'b0),                                          //           (terminated)
		.locked             (),                                              //           (terminated)
		.phasedone          (),                                              //           (terminated)
		.phasecounterselect (4'b0000),                                       //           (terminated)
		.phaseupdown        (1'b0),                                          //           (terminated)
		.phasestep          (1'b0),                                          //           (terminated)
		.scanclk            (1'b0),                                          //           (terminated)
		.scanclkena         (1'b0),                                          //           (terminated)
		.scandata           (1'b0),                                          //           (terminated)
		.configupdate       (1'b0)                                           //           (terminated)
	);

	ECE385_io_hex io_hex (
		.clk        (nios2_pll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_io_hex_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_hex_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_hex_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_hex_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_hex_s1_readdata),   //                    .readdata
		.out_port   (io_hex_export)                           // external_connection.export
	);

	ECE385_io_keys io_keys (
		.clk      (nios2_pll_c0_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_io_keys_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_io_keys_s1_readdata), //                    .readdata
		.in_port  (io_keys_export)                         // external_connection.export
	);

	ECE385_io_led_green io_led_green (
		.clk        (nios2_pll_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_io_led_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_led_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_led_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_led_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_led_green_s1_readdata),   //                    .readdata
		.out_port   (io_led_green_export)                           // external_connection.export
	);

	ECE385_io_led_red io_led_red (
		.clk        (nios2_pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_io_led_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_led_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_led_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_led_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_led_red_s1_readdata),   //                    .readdata
		.out_port   (io_led_red_export)                           // external_connection.export
	);

	ECE385_io_switches io_switches (
		.clk      (nios2_pll_c0_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_io_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_io_switches_s1_readdata), //                    .readdata
		.in_port  (io_switches_export)                         // external_connection.export
	);

	ECE385_keycode keycode (
		.clk        (nios2_pll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	ECE385_nios2_cpu nios2_cpu (
		.clk                                 (nios2_pll_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	ECE385_nios2_jtag_uart nios2_jtag_uart (
		.clk            (nios2_pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                 //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                         //               irq.irq
	);

	ECE385_nios2_onchip_mem nios2_onchip_mem (
		.clk        (nios2_pll_c0_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_nios2_onchip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_nios2_onchip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_nios2_onchip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_nios2_onchip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_nios2_onchip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_nios2_onchip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_nios2_onchip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	ECE385_nios2_pll nios2_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read               (mm_interconnect_0_nios2_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_nios2_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_nios2_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_nios2_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_nios2_pll_pll_slave_writedata), //                      .writedata
		.inclk0             (clk_clk),                                         //                inclk0.clk
		.c0                 (nios2_pll_c0_clk),                                //                    c0.clk
		.c1                 (nios2_pll_sdram_clk),                             //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (4'b0000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	ECE385_nios2_sysid nios2_sysid (
		.clock    (nios2_pll_c0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //         reset.reset_n
		.readdata (mm_interconnect_0_nios2_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_nios2_sysid_control_slave_address)   //              .address
	);

	ECE385_nios2_timer nios2_timer (
		.clk        (nios2_pll_c0_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             // reset.reset_n
		.address    (mm_interconnect_0_nios2_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_nios2_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_nios2_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_nios2_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_nios2_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                     //   irq.irq
	);

	ECE385_otg_hpi_address otg_hpi_address (
		.clk        (nios2_pll_c0_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	ECE385_otg_hpi_cs otg_hpi_cs (
		.clk        (nios2_pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	ECE385_otg_hpi_data otg_hpi_data (
		.clk        (nios2_pll_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	ECE385_otg_hpi_cs otg_hpi_r (
		.clk        (nios2_pll_c0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	ECE385_otg_hpi_cs otg_hpi_reset (
		.clk        (nios2_pll_c0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	ECE385_otg_hpi_cs otg_hpi_w (
		.clk        (nios2_pll_c0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	ECE385_sdram sdram (
		.clk            (nios2_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	ECE385_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                               (clk_clk),                                                         //                                             clk_0_clk.clk
		.nios2_pll_c0_clk                                            (nios2_pll_c0_clk),                                                //                                          nios2_pll_c0.clk
		.nios2_cpu_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                              //                 nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_jtag_uart_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                  //           nios2_jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                              // nios2_pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                               (nios2_cpu_data_master_address),                                   //                                 nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest                           (nios2_cpu_data_master_waitrequest),                               //                                                      .waitrequest
		.nios2_cpu_data_master_byteenable                            (nios2_cpu_data_master_byteenable),                                //                                                      .byteenable
		.nios2_cpu_data_master_read                                  (nios2_cpu_data_master_read),                                      //                                                      .read
		.nios2_cpu_data_master_readdata                              (nios2_cpu_data_master_readdata),                                  //                                                      .readdata
		.nios2_cpu_data_master_write                                 (nios2_cpu_data_master_write),                                     //                                                      .write
		.nios2_cpu_data_master_writedata                             (nios2_cpu_data_master_writedata),                                 //                                                      .writedata
		.nios2_cpu_data_master_debugaccess                           (nios2_cpu_data_master_debugaccess),                               //                                                      .debugaccess
		.nios2_cpu_instruction_master_address                        (nios2_cpu_instruction_master_address),                            //                          nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest                    (nios2_cpu_instruction_master_waitrequest),                        //                                                      .waitrequest
		.nios2_cpu_instruction_master_read                           (nios2_cpu_instruction_master_read),                               //                                                      .read
		.nios2_cpu_instruction_master_readdata                       (nios2_cpu_instruction_master_readdata),                           //                                                      .readdata
		.eth0_mdio_avalon_slave_address                              (mm_interconnect_0_eth0_mdio_avalon_slave_address),                //                                eth0_mdio_avalon_slave.address
		.eth0_mdio_avalon_slave_write                                (mm_interconnect_0_eth0_mdio_avalon_slave_write),                  //                                                      .write
		.eth0_mdio_avalon_slave_read                                 (mm_interconnect_0_eth0_mdio_avalon_slave_read),                   //                                                      .read
		.eth0_mdio_avalon_slave_readdata                             (mm_interconnect_0_eth0_mdio_avalon_slave_readdata),               //                                                      .readdata
		.eth0_mdio_avalon_slave_writedata                            (mm_interconnect_0_eth0_mdio_avalon_slave_writedata),              //                                                      .writedata
		.eth0_mdio_avalon_slave_waitrequest                          (mm_interconnect_0_eth0_mdio_avalon_slave_waitrequest),            //                                                      .waitrequest
		.eth1_mdio_avalon_slave_address                              (mm_interconnect_0_eth1_mdio_avalon_slave_address),                //                                eth1_mdio_avalon_slave.address
		.eth1_mdio_avalon_slave_write                                (mm_interconnect_0_eth1_mdio_avalon_slave_write),                  //                                                      .write
		.eth1_mdio_avalon_slave_read                                 (mm_interconnect_0_eth1_mdio_avalon_slave_read),                   //                                                      .read
		.eth1_mdio_avalon_slave_readdata                             (mm_interconnect_0_eth1_mdio_avalon_slave_readdata),               //                                                      .readdata
		.eth1_mdio_avalon_slave_writedata                            (mm_interconnect_0_eth1_mdio_avalon_slave_writedata),              //                                                      .writedata
		.eth1_mdio_avalon_slave_waitrequest                          (mm_interconnect_0_eth1_mdio_avalon_slave_waitrequest),            //                                                      .waitrequest
		.eth_pll_pll_slave_address                                   (mm_interconnect_0_eth_pll_pll_slave_address),                     //                                     eth_pll_pll_slave.address
		.eth_pll_pll_slave_write                                     (mm_interconnect_0_eth_pll_pll_slave_write),                       //                                                      .write
		.eth_pll_pll_slave_read                                      (mm_interconnect_0_eth_pll_pll_slave_read),                        //                                                      .read
		.eth_pll_pll_slave_readdata                                  (mm_interconnect_0_eth_pll_pll_slave_readdata),                    //                                                      .readdata
		.eth_pll_pll_slave_writedata                                 (mm_interconnect_0_eth_pll_pll_slave_writedata),                   //                                                      .writedata
		.io_hex_s1_address                                           (mm_interconnect_0_io_hex_s1_address),                             //                                             io_hex_s1.address
		.io_hex_s1_write                                             (mm_interconnect_0_io_hex_s1_write),                               //                                                      .write
		.io_hex_s1_readdata                                          (mm_interconnect_0_io_hex_s1_readdata),                            //                                                      .readdata
		.io_hex_s1_writedata                                         (mm_interconnect_0_io_hex_s1_writedata),                           //                                                      .writedata
		.io_hex_s1_chipselect                                        (mm_interconnect_0_io_hex_s1_chipselect),                          //                                                      .chipselect
		.io_keys_s1_address                                          (mm_interconnect_0_io_keys_s1_address),                            //                                            io_keys_s1.address
		.io_keys_s1_readdata                                         (mm_interconnect_0_io_keys_s1_readdata),                           //                                                      .readdata
		.io_led_green_s1_address                                     (mm_interconnect_0_io_led_green_s1_address),                       //                                       io_led_green_s1.address
		.io_led_green_s1_write                                       (mm_interconnect_0_io_led_green_s1_write),                         //                                                      .write
		.io_led_green_s1_readdata                                    (mm_interconnect_0_io_led_green_s1_readdata),                      //                                                      .readdata
		.io_led_green_s1_writedata                                   (mm_interconnect_0_io_led_green_s1_writedata),                     //                                                      .writedata
		.io_led_green_s1_chipselect                                  (mm_interconnect_0_io_led_green_s1_chipselect),                    //                                                      .chipselect
		.io_led_red_s1_address                                       (mm_interconnect_0_io_led_red_s1_address),                         //                                         io_led_red_s1.address
		.io_led_red_s1_write                                         (mm_interconnect_0_io_led_red_s1_write),                           //                                                      .write
		.io_led_red_s1_readdata                                      (mm_interconnect_0_io_led_red_s1_readdata),                        //                                                      .readdata
		.io_led_red_s1_writedata                                     (mm_interconnect_0_io_led_red_s1_writedata),                       //                                                      .writedata
		.io_led_red_s1_chipselect                                    (mm_interconnect_0_io_led_red_s1_chipselect),                      //                                                      .chipselect
		.io_switches_s1_address                                      (mm_interconnect_0_io_switches_s1_address),                        //                                        io_switches_s1.address
		.io_switches_s1_readdata                                     (mm_interconnect_0_io_switches_s1_readdata),                       //                                                      .readdata
		.keycode_s1_address                                          (mm_interconnect_0_keycode_s1_address),                            //                                            keycode_s1.address
		.keycode_s1_write                                            (mm_interconnect_0_keycode_s1_write),                              //                                                      .write
		.keycode_s1_readdata                                         (mm_interconnect_0_keycode_s1_readdata),                           //                                                      .readdata
		.keycode_s1_writedata                                        (mm_interconnect_0_keycode_s1_writedata),                          //                                                      .writedata
		.keycode_s1_chipselect                                       (mm_interconnect_0_keycode_s1_chipselect),                         //                                                      .chipselect
		.nios2_cpu_debug_mem_slave_address                           (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),             //                             nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write                             (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),               //                                                      .write
		.nios2_cpu_debug_mem_slave_read                              (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),                //                                                      .read
		.nios2_cpu_debug_mem_slave_readdata                          (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),            //                                                      .readdata
		.nios2_cpu_debug_mem_slave_writedata                         (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),           //                                                      .writedata
		.nios2_cpu_debug_mem_slave_byteenable                        (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),          //                                                      .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),         //                                                      .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),         //                                                      .debugaccess
		.nios2_jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_address),     //                     nios2_jtag_uart_avalon_jtag_slave.address
		.nios2_jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_write),       //                                                      .write
		.nios2_jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_read),        //                                                      .read
		.nios2_jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_readdata),    //                                                      .readdata
		.nios2_jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_writedata),   //                                                      .writedata
		.nios2_jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_waitrequest), //                                                      .waitrequest
		.nios2_jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_chipselect),  //                                                      .chipselect
		.nios2_onchip_mem_s1_address                                 (mm_interconnect_0_nios2_onchip_mem_s1_address),                   //                                   nios2_onchip_mem_s1.address
		.nios2_onchip_mem_s1_write                                   (mm_interconnect_0_nios2_onchip_mem_s1_write),                     //                                                      .write
		.nios2_onchip_mem_s1_readdata                                (mm_interconnect_0_nios2_onchip_mem_s1_readdata),                  //                                                      .readdata
		.nios2_onchip_mem_s1_writedata                               (mm_interconnect_0_nios2_onchip_mem_s1_writedata),                 //                                                      .writedata
		.nios2_onchip_mem_s1_byteenable                              (mm_interconnect_0_nios2_onchip_mem_s1_byteenable),                //                                                      .byteenable
		.nios2_onchip_mem_s1_chipselect                              (mm_interconnect_0_nios2_onchip_mem_s1_chipselect),                //                                                      .chipselect
		.nios2_onchip_mem_s1_clken                                   (mm_interconnect_0_nios2_onchip_mem_s1_clken),                     //                                                      .clken
		.nios2_pll_pll_slave_address                                 (mm_interconnect_0_nios2_pll_pll_slave_address),                   //                                   nios2_pll_pll_slave.address
		.nios2_pll_pll_slave_write                                   (mm_interconnect_0_nios2_pll_pll_slave_write),                     //                                                      .write
		.nios2_pll_pll_slave_read                                    (mm_interconnect_0_nios2_pll_pll_slave_read),                      //                                                      .read
		.nios2_pll_pll_slave_readdata                                (mm_interconnect_0_nios2_pll_pll_slave_readdata),                  //                                                      .readdata
		.nios2_pll_pll_slave_writedata                               (mm_interconnect_0_nios2_pll_pll_slave_writedata),                 //                                                      .writedata
		.nios2_sysid_control_slave_address                           (mm_interconnect_0_nios2_sysid_control_slave_address),             //                             nios2_sysid_control_slave.address
		.nios2_sysid_control_slave_readdata                          (mm_interconnect_0_nios2_sysid_control_slave_readdata),            //                                                      .readdata
		.nios2_timer_s1_address                                      (mm_interconnect_0_nios2_timer_s1_address),                        //                                        nios2_timer_s1.address
		.nios2_timer_s1_write                                        (mm_interconnect_0_nios2_timer_s1_write),                          //                                                      .write
		.nios2_timer_s1_readdata                                     (mm_interconnect_0_nios2_timer_s1_readdata),                       //                                                      .readdata
		.nios2_timer_s1_writedata                                    (mm_interconnect_0_nios2_timer_s1_writedata),                      //                                                      .writedata
		.nios2_timer_s1_chipselect                                   (mm_interconnect_0_nios2_timer_s1_chipselect),                     //                                                      .chipselect
		.otg_hpi_address_s1_address                                  (mm_interconnect_0_otg_hpi_address_s1_address),                    //                                    otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                                    (mm_interconnect_0_otg_hpi_address_s1_write),                      //                                                      .write
		.otg_hpi_address_s1_readdata                                 (mm_interconnect_0_otg_hpi_address_s1_readdata),                   //                                                      .readdata
		.otg_hpi_address_s1_writedata                                (mm_interconnect_0_otg_hpi_address_s1_writedata),                  //                                                      .writedata
		.otg_hpi_address_s1_chipselect                               (mm_interconnect_0_otg_hpi_address_s1_chipselect),                 //                                                      .chipselect
		.otg_hpi_cs_s1_address                                       (mm_interconnect_0_otg_hpi_cs_s1_address),                         //                                         otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                                         (mm_interconnect_0_otg_hpi_cs_s1_write),                           //                                                      .write
		.otg_hpi_cs_s1_readdata                                      (mm_interconnect_0_otg_hpi_cs_s1_readdata),                        //                                                      .readdata
		.otg_hpi_cs_s1_writedata                                     (mm_interconnect_0_otg_hpi_cs_s1_writedata),                       //                                                      .writedata
		.otg_hpi_cs_s1_chipselect                                    (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                      //                                                      .chipselect
		.otg_hpi_data_s1_address                                     (mm_interconnect_0_otg_hpi_data_s1_address),                       //                                       otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                                       (mm_interconnect_0_otg_hpi_data_s1_write),                         //                                                      .write
		.otg_hpi_data_s1_readdata                                    (mm_interconnect_0_otg_hpi_data_s1_readdata),                      //                                                      .readdata
		.otg_hpi_data_s1_writedata                                   (mm_interconnect_0_otg_hpi_data_s1_writedata),                     //                                                      .writedata
		.otg_hpi_data_s1_chipselect                                  (mm_interconnect_0_otg_hpi_data_s1_chipselect),                    //                                                      .chipselect
		.otg_hpi_r_s1_address                                        (mm_interconnect_0_otg_hpi_r_s1_address),                          //                                          otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                                          (mm_interconnect_0_otg_hpi_r_s1_write),                            //                                                      .write
		.otg_hpi_r_s1_readdata                                       (mm_interconnect_0_otg_hpi_r_s1_readdata),                         //                                                      .readdata
		.otg_hpi_r_s1_writedata                                      (mm_interconnect_0_otg_hpi_r_s1_writedata),                        //                                                      .writedata
		.otg_hpi_r_s1_chipselect                                     (mm_interconnect_0_otg_hpi_r_s1_chipselect),                       //                                                      .chipselect
		.otg_hpi_reset_s1_address                                    (mm_interconnect_0_otg_hpi_reset_s1_address),                      //                                      otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                                      (mm_interconnect_0_otg_hpi_reset_s1_write),                        //                                                      .write
		.otg_hpi_reset_s1_readdata                                   (mm_interconnect_0_otg_hpi_reset_s1_readdata),                     //                                                      .readdata
		.otg_hpi_reset_s1_writedata                                  (mm_interconnect_0_otg_hpi_reset_s1_writedata),                    //                                                      .writedata
		.otg_hpi_reset_s1_chipselect                                 (mm_interconnect_0_otg_hpi_reset_s1_chipselect),                   //                                                      .chipselect
		.otg_hpi_w_s1_address                                        (mm_interconnect_0_otg_hpi_w_s1_address),                          //                                          otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                                          (mm_interconnect_0_otg_hpi_w_s1_write),                            //                                                      .write
		.otg_hpi_w_s1_readdata                                       (mm_interconnect_0_otg_hpi_w_s1_readdata),                         //                                                      .readdata
		.otg_hpi_w_s1_writedata                                      (mm_interconnect_0_otg_hpi_w_s1_writedata),                        //                                                      .writedata
		.otg_hpi_w_s1_chipselect                                     (mm_interconnect_0_otg_hpi_w_s1_chipselect),                       //                                                      .chipselect
		.sdram_s1_address                                            (mm_interconnect_0_sdram_s1_address),                              //                                              sdram_s1.address
		.sdram_s1_write                                              (mm_interconnect_0_sdram_s1_write),                                //                                                      .write
		.sdram_s1_read                                               (mm_interconnect_0_sdram_s1_read),                                 //                                                      .read
		.sdram_s1_readdata                                           (mm_interconnect_0_sdram_s1_readdata),                             //                                                      .readdata
		.sdram_s1_writedata                                          (mm_interconnect_0_sdram_s1_writedata),                            //                                                      .writedata
		.sdram_s1_byteenable                                         (mm_interconnect_0_sdram_s1_byteenable),                           //                                                      .byteenable
		.sdram_s1_readdatavalid                                      (mm_interconnect_0_sdram_s1_readdatavalid),                        //                                                      .readdatavalid
		.sdram_s1_waitrequest                                        (mm_interconnect_0_sdram_s1_waitrequest),                          //                                                      .waitrequest
		.sdram_s1_chipselect                                         (mm_interconnect_0_sdram_s1_chipselect)                            //                                                      .chipselect
	);

	ECE385_irq_mapper irq_mapper (
		.clk           (nios2_pll_c0_clk),                   //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_cpu_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (nios2_pll_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset),    // reset_in1.reset
		.clk            (nios2_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
