// ECE385.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ECE385 (
		input  wire        audio_mem_clk2_clk,                             //                          audio_mem_clk2.clk
		input  wire        audio_mem_reset2_reset,                         //                        audio_mem_reset2.reset
		input  wire [11:0] audio_mem_s2_address,                           //                            audio_mem_s2.address
		input  wire        audio_mem_s2_chipselect,                        //                                        .chipselect
		input  wire        audio_mem_s2_clken,                             //                                        .clken
		input  wire        audio_mem_s2_write,                             //                                        .write
		output wire [31:0] audio_mem_s2_readdata,                          //                                        .readdata
		input  wire [31:0] audio_mem_s2_writedata,                         //                                        .writedata
		input  wire [3:0]  audio_mem_s2_byteenable,                        //                                        .byteenable
		input  wire [31:0] audio_position_export,                          //                          audio_position.export
		output wire [31:0] audio_position_end_export,                      //                      audio_position_end.export
		input  wire        clk_clk,                                        //                                     clk.clk
		output wire        eth0_mdio_mdc,                                  //                               eth0_mdio.mdc
		input  wire        eth0_mdio_mdio_in,                              //                                        .mdio_in
		output wire        eth0_mdio_mdio_out,                             //                                        .mdio_out
		output wire        eth0_mdio_mdio_oen,                             //                                        .mdio_oen
		input  wire [4:0]  eth0_mdio_phy_addr,                             //                                        .phy_addr
		input  wire [7:0]  eth0_rx_fifo_in_data,                           //                         eth0_rx_fifo_in.data
		input  wire        eth0_rx_fifo_in_valid,                          //                                        .valid
		output wire        eth0_rx_fifo_in_ready,                          //                                        .ready
		input  wire        eth0_rx_fifo_in_startofpacket,                  //                                        .startofpacket
		input  wire        eth0_rx_fifo_in_endofpacket,                    //                                        .endofpacket
		input  wire [2:0]  eth0_rx_fifo_in_error,                          //                                        .error
		input  wire        eth0_rx_fifo_in_clk_clk,                        //                     eth0_rx_fifo_in_clk.clk
		input  wire        eth0_rx_fifo_in_clk_reset_reset_n,              //               eth0_rx_fifo_in_clk_reset.reset_n
		input  wire [31:0] eth0_tx_dma_buffer_in_0_data,                   //                 eth0_tx_dma_buffer_in_0.data
		input  wire        eth0_tx_dma_buffer_in_0_valid,                  //                                        .valid
		output wire        eth0_tx_dma_buffer_in_0_ready,                  //                                        .ready
		input  wire        eth0_tx_dma_buffer_in_0_startofpacket,          //                                        .startofpacket
		input  wire        eth0_tx_dma_buffer_in_0_endofpacket,            //                                        .endofpacket
		input  wire [1:0]  eth0_tx_dma_buffer_in_0_empty,                  //                                        .empty
		input  wire        eth0_tx_dma_buffer_in_clk_0_clk,                //             eth0_tx_dma_buffer_in_clk_0.clk
		input  wire        eth0_tx_dma_buffer_in_rst_0_reset,              //             eth0_tx_dma_buffer_in_rst_0.reset
		output wire [7:0]  eth0_tx_dma_buffer_out_0_data,                  //                eth0_tx_dma_buffer_out_0.data
		output wire        eth0_tx_dma_buffer_out_0_valid,                 //                                        .valid
		input  wire        eth0_tx_dma_buffer_out_0_ready,                 //                                        .ready
		output wire        eth0_tx_dma_buffer_out_0_startofpacket,         //                                        .startofpacket
		output wire        eth0_tx_dma_buffer_out_0_endofpacket,           //                                        .endofpacket
		output wire [31:0] eth0_tx_fifo_out_data,                          //                        eth0_tx_fifo_out.data
		output wire        eth0_tx_fifo_out_valid,                         //                                        .valid
		input  wire        eth0_tx_fifo_out_ready,                         //                                        .ready
		output wire        eth0_tx_fifo_out_startofpacket,                 //                                        .startofpacket
		output wire        eth0_tx_fifo_out_endofpacket,                   //                                        .endofpacket
		output wire [1:0]  eth0_tx_fifo_out_empty,                         //                                        .empty
		input  wire        eth0_tx_fifo_out_clk_clk,                       //                    eth0_tx_fifo_out_clk.clk
		input  wire        eth0_tx_fifo_out_clk_reset_reset_n,             //              eth0_tx_fifo_out_clk_reset.reset_n
		output wire        eth1_mdio_mdc,                                  //                               eth1_mdio.mdc
		input  wire        eth1_mdio_mdio_in,                              //                                        .mdio_in
		output wire        eth1_mdio_mdio_out,                             //                                        .mdio_out
		output wire        eth1_mdio_mdio_oen,                             //                                        .mdio_oen
		input  wire [4:0]  eth1_mdio_phy_addr,                             //                                        .phy_addr
		input  wire [7:0]  eth1_rx_fifo_in_data,                           //                         eth1_rx_fifo_in.data
		input  wire        eth1_rx_fifo_in_valid,                          //                                        .valid
		output wire        eth1_rx_fifo_in_ready,                          //                                        .ready
		input  wire        eth1_rx_fifo_in_startofpacket,                  //                                        .startofpacket
		input  wire        eth1_rx_fifo_in_endofpacket,                    //                                        .endofpacket
		input  wire [2:0]  eth1_rx_fifo_in_error,                          //                                        .error
		input  wire        eth1_rx_fifo_in_clk_clk,                        //                     eth1_rx_fifo_in_clk.clk
		input  wire        eth1_rx_fifo_in_clk_reset_reset_n,              //               eth1_rx_fifo_in_clk_reset.reset_n
		input  wire [31:0] eth1_tx_dma_buffer_in_0_data,                   //                 eth1_tx_dma_buffer_in_0.data
		input  wire        eth1_tx_dma_buffer_in_0_valid,                  //                                        .valid
		output wire        eth1_tx_dma_buffer_in_0_ready,                  //                                        .ready
		input  wire        eth1_tx_dma_buffer_in_0_startofpacket,          //                                        .startofpacket
		input  wire        eth1_tx_dma_buffer_in_0_endofpacket,            //                                        .endofpacket
		input  wire [1:0]  eth1_tx_dma_buffer_in_0_empty,                  //                                        .empty
		input  wire        eth1_tx_dma_buffer_in_clk_0_clk,                //             eth1_tx_dma_buffer_in_clk_0.clk
		input  wire        eth1_tx_dma_buffer_in_rst_0_reset,              //             eth1_tx_dma_buffer_in_rst_0.reset
		output wire [7:0]  eth1_tx_dma_buffer_out_0_data,                  //                eth1_tx_dma_buffer_out_0.data
		output wire        eth1_tx_dma_buffer_out_0_valid,                 //                                        .valid
		input  wire        eth1_tx_dma_buffer_out_0_ready,                 //                                        .ready
		output wire        eth1_tx_dma_buffer_out_0_startofpacket,         //                                        .startofpacket
		output wire        eth1_tx_dma_buffer_out_0_endofpacket,           //                                        .endofpacket
		output wire [31:0] eth1_tx_fifo_out_data,                          //                        eth1_tx_fifo_out.data
		output wire        eth1_tx_fifo_out_valid,                         //                                        .valid
		input  wire        eth1_tx_fifo_out_ready,                         //                                        .ready
		output wire        eth1_tx_fifo_out_startofpacket,                 //                                        .startofpacket
		output wire        eth1_tx_fifo_out_endofpacket,                   //                                        .endofpacket
		output wire [1:0]  eth1_tx_fifo_out_empty,                         //                                        .empty
		input  wire        eth1_tx_fifo_out_clk_clk,                       //                    eth1_tx_fifo_out_clk.clk
		input  wire        eth1_tx_fifo_out_clk_reset_reset_n,             //              eth1_tx_fifo_out_clk_reset.reset_n
		output wire [31:0] io_hex_export,                                  //                                  io_hex.export
		input  wire [3:0]  io_keys_export,                                 //                                 io_keys.export
		output wire [8:0]  io_led_green_export,                            //                            io_led_green.export
		output wire [17:0] io_led_red_export,                              //                              io_led_red.export
		input  wire [17:0] io_switches_export,                             //                             io_switches.export
		input  wire        io_vga_sync_export,                             //                             io_vga_sync.export
		output wire        nios2_pll_ethernet_clk,                         //                      nios2_pll_ethernet.clk
		output wire        nios2_pll_sdram_clk,                            //                         nios2_pll_sdram.clk
		output wire        nios2_pll_vga_clk,                              //                           nios2_pll_vga.clk
		output wire [1:0]  otg_hpi_address_export,                         //                         otg_hpi_address.export
		output wire        otg_hpi_cs_export,                              //                              otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,                           //                            otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,                          //                                        .out_port
		output wire        otg_hpi_r_export,                               //                               otg_hpi_r.export
		output wire        otg_hpi_reset_export,                           //                           otg_hpi_reset.export
		output wire        otg_hpi_w_export,                               //                               otg_hpi_w.export
		input  wire        reset_reset_n,                                  //                                   reset.reset_n
		output wire [12:0] sdram_addr,                                     //                                   sdram.addr
		output wire [1:0]  sdram_ba,                                       //                                        .ba
		output wire        sdram_cas_n,                                    //                                        .cas_n
		output wire        sdram_cke,                                      //                                        .cke
		output wire        sdram_cs_n,                                     //                                        .cs_n
		inout  wire [31:0] sdram_dq,                                       //                                        .dq
		output wire [3:0]  sdram_dqm,                                      //                                        .dqm
		output wire        sdram_ras_n,                                    //                                        .ras_n
		output wire        sdram_we_n,                                     //                                        .we_n
		output wire [19:0] sram_sram_addr,                                 //                                    sram.sram_addr
		output wire        sram_sram_ce_n,                                 //                                        .sram_ce_n
		inout  wire [15:0] sram_sram_dq,                                   //                                        .sram_dq
		output wire        sram_sram_lb_n,                                 //                                        .sram_lb_n
		output wire        sram_sram_oe_n,                                 //                                        .sram_oe_n
		output wire        sram_sram_ub_n,                                 //                                        .sram_ub_n
		output wire        sram_sram_we_n,                                 //                                        .sram_we_n
		input  wire        usb_clk_clk,                                    //                                 usb_clk.clk
		output wire        usb_nios2_cpu_custom_instruction_master_readra, // usb_nios2_cpu_custom_instruction_master.readra
		input  wire        usb_reset_reset_n,                              //                               usb_reset.reset_n
		input  wire [9:0]  vga_vga_drawx,                                  //                                     vga.vga_drawx
		input  wire [9:0]  vga_vga_drawy,                                  //                                        .vga_drawy
		output wire [15:0] vga_vga_val,                                    //                                        .vga_val
		output wire [31:0] vga_background_offset_export,                   //                   vga_background_offset.export
		input  wire        vga_sprite_0_clk2_clk,                          //                       vga_sprite_0_clk2.clk
		input  wire        vga_sprite_0_reset2_reset,                      //                     vga_sprite_0_reset2.reset
		input  wire [10:0] vga_sprite_0_s2_address,                        //                         vga_sprite_0_s2.address
		input  wire        vga_sprite_0_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_0_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_0_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_0_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_0_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_0_s2_byteenable,                     //                                        .byteenable
		input  wire        vga_sprite_1_clk2_clk,                          //                       vga_sprite_1_clk2.clk
		input  wire        vga_sprite_1_reset2_reset,                      //                     vga_sprite_1_reset2.reset
		input  wire [10:0] vga_sprite_1_s2_address,                        //                         vga_sprite_1_s2.address
		input  wire        vga_sprite_1_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_1_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_1_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_1_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_1_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_1_s2_byteenable,                     //                                        .byteenable
		input  wire        vga_sprite_2_clk2_clk,                          //                       vga_sprite_2_clk2.clk
		input  wire        vga_sprite_2_reset2_reset,                      //                     vga_sprite_2_reset2.reset
		input  wire [10:0] vga_sprite_2_s2_address,                        //                         vga_sprite_2_s2.address
		input  wire        vga_sprite_2_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_2_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_2_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_2_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_2_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_2_s2_byteenable,                     //                                        .byteenable
		input  wire        vga_sprite_3_clk2_clk,                          //                       vga_sprite_3_clk2.clk
		input  wire        vga_sprite_3_reset2_reset,                      //                     vga_sprite_3_reset2.reset
		input  wire [10:0] vga_sprite_3_s2_address,                        //                         vga_sprite_3_s2.address
		input  wire        vga_sprite_3_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_3_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_3_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_3_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_3_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_3_s2_byteenable,                     //                                        .byteenable
		input  wire        vga_sprite_4_clk2_clk,                          //                       vga_sprite_4_clk2.clk
		input  wire        vga_sprite_4_reset2_reset,                      //                     vga_sprite_4_reset2.reset
		input  wire [10:0] vga_sprite_4_s2_address,                        //                         vga_sprite_4_s2.address
		input  wire        vga_sprite_4_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_4_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_4_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_4_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_4_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_4_s2_byteenable,                     //                                        .byteenable
		input  wire        vga_sprite_5_clk2_clk,                          //                       vga_sprite_5_clk2.clk
		input  wire        vga_sprite_5_reset2_reset,                      //                     vga_sprite_5_reset2.reset
		input  wire [10:0] vga_sprite_5_s2_address,                        //                         vga_sprite_5_s2.address
		input  wire        vga_sprite_5_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_5_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_5_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_5_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_5_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_5_s2_byteenable,                     //                                        .byteenable
		input  wire        vga_sprite_6_clk2_clk,                          //                       vga_sprite_6_clk2.clk
		input  wire        vga_sprite_6_reset2_reset,                      //                     vga_sprite_6_reset2.reset
		input  wire [10:0] vga_sprite_6_s2_address,                        //                         vga_sprite_6_s2.address
		input  wire        vga_sprite_6_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_6_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_6_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_6_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_6_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_6_s2_byteenable,                     //                                        .byteenable
		input  wire        vga_sprite_7_clk2_clk,                          //                       vga_sprite_7_clk2.clk
		input  wire        vga_sprite_7_reset2_reset,                      //                     vga_sprite_7_reset2.reset
		input  wire [10:0] vga_sprite_7_s2_address,                        //                         vga_sprite_7_s2.address
		input  wire        vga_sprite_7_s2_chipselect,                     //                                        .chipselect
		input  wire        vga_sprite_7_s2_clken,                          //                                        .clken
		input  wire        vga_sprite_7_s2_write,                          //                                        .write
		output wire [15:0] vga_sprite_7_s2_readdata,                       //                                        .readdata
		input  wire [15:0] vga_sprite_7_s2_writedata,                      //                                        .writedata
		input  wire [1:0]  vga_sprite_7_s2_byteenable,                     //                                        .byteenable
		output wire [7:0]  vga_sprite_params_pass_address,                 //                  vga_sprite_params_pass.address
		output wire        vga_sprite_params_pass_read,                    //                                        .read
		input  wire [31:0] vga_sprite_params_pass_readdata,                //                                        .readdata
		output wire        vga_sprite_params_pass_write,                   //                                        .write
		output wire [31:0] vga_sprite_params_pass_writedata,               //                                        .writedata
		output wire        vga_sprite_params_reset_reset                   //                 vga_sprite_params_reset.reset
	);

	wire         eth0_rx_fifo_out_valid;                                          // eth0_rx_fifo:out_valid -> eth0_rx_dma:in_valid
	wire   [7:0] eth0_rx_fifo_out_data;                                           // eth0_rx_fifo:out_data -> eth0_rx_dma:in_data
	wire         eth0_rx_fifo_out_ready;                                          // eth0_rx_dma:in_ready -> eth0_rx_fifo:out_ready
	wire         eth0_rx_fifo_out_startofpacket;                                  // eth0_rx_fifo:out_startofpacket -> eth0_rx_dma:in_startofpacket
	wire         eth0_rx_fifo_out_endofpacket;                                    // eth0_rx_fifo:out_endofpacket -> eth0_rx_dma:in_endofpacket
	wire   [2:0] eth0_rx_fifo_out_error;                                          // eth0_rx_fifo:out_error -> eth0_rx_dma:in_error
	wire         eth0_tx_dma_out_valid;                                           // eth0_tx_dma:out_valid -> eth0_tx_fifo:in_valid
	wire  [31:0] eth0_tx_dma_out_data;                                            // eth0_tx_dma:out_data -> eth0_tx_fifo:in_data
	wire         eth0_tx_dma_out_ready;                                           // eth0_tx_fifo:in_ready -> eth0_tx_dma:out_ready
	wire         eth0_tx_dma_out_startofpacket;                                   // eth0_tx_dma:out_startofpacket -> eth0_tx_fifo:in_startofpacket
	wire         eth0_tx_dma_out_endofpacket;                                     // eth0_tx_dma:out_endofpacket -> eth0_tx_fifo:in_endofpacket
	wire   [1:0] eth0_tx_dma_out_empty;                                           // eth0_tx_dma:out_empty -> eth0_tx_fifo:in_empty
	wire         eth1_rx_fifo_out_valid;                                          // eth1_rx_fifo:out_valid -> eth1_rx_dma:in_valid
	wire   [7:0] eth1_rx_fifo_out_data;                                           // eth1_rx_fifo:out_data -> eth1_rx_dma:in_data
	wire         eth1_rx_fifo_out_ready;                                          // eth1_rx_dma:in_ready -> eth1_rx_fifo:out_ready
	wire         eth1_rx_fifo_out_startofpacket;                                  // eth1_rx_fifo:out_startofpacket -> eth1_rx_dma:in_startofpacket
	wire         eth1_rx_fifo_out_endofpacket;                                    // eth1_rx_fifo:out_endofpacket -> eth1_rx_dma:in_endofpacket
	wire   [2:0] eth1_rx_fifo_out_error;                                          // eth1_rx_fifo:out_error -> eth1_rx_dma:in_error
	wire         eth1_tx_dma_out_valid;                                           // eth1_tx_dma:out_valid -> eth1_tx_fifo:in_valid
	wire  [31:0] eth1_tx_dma_out_data;                                            // eth1_tx_dma:out_data -> eth1_tx_fifo:in_data
	wire         eth1_tx_dma_out_ready;                                           // eth1_tx_fifo:in_ready -> eth1_tx_dma:out_ready
	wire         eth1_tx_dma_out_startofpacket;                                   // eth1_tx_dma:out_startofpacket -> eth1_tx_fifo:in_startofpacket
	wire         eth1_tx_dma_out_endofpacket;                                     // eth1_tx_dma:out_endofpacket -> eth1_tx_fifo:in_endofpacket
	wire   [1:0] eth1_tx_dma_out_empty;                                           // eth1_tx_dma:out_empty -> eth1_tx_fifo:in_empty
	wire         nios2_pll_c2_clk;                                                // nios2_pll:c2 -> sram_multiplexer:CLK2
	wire  [31:0] nios2_cpu_data_master_readdata;                                  // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                               // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                               // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [27:0] nios2_cpu_data_master_address;                                   // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                                // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                      // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_write;                                     // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                 // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_dma_m_read_readdata;                                       // mm_interconnect_0:nios2_dma_m_read_readdata -> nios2_dma:m_read_readdata
	wire         nios2_dma_m_read_waitrequest;                                    // mm_interconnect_0:nios2_dma_m_read_waitrequest -> nios2_dma:m_read_waitrequest
	wire  [31:0] nios2_dma_m_read_address;                                        // nios2_dma:m_read_address -> mm_interconnect_0:nios2_dma_m_read_address
	wire         nios2_dma_m_read_read;                                           // nios2_dma:m_read_read -> mm_interconnect_0:nios2_dma_m_read_read
	wire         nios2_dma_m_read_readdatavalid;                                  // mm_interconnect_0:nios2_dma_m_read_readdatavalid -> nios2_dma:m_read_readdatavalid
	wire         nios2_dma_m_write_waitrequest;                                   // mm_interconnect_0:nios2_dma_m_write_waitrequest -> nios2_dma:m_write_waitrequest
	wire  [31:0] nios2_dma_m_write_address;                                       // nios2_dma:m_write_address -> mm_interconnect_0:nios2_dma_m_write_address
	wire   [3:0] nios2_dma_m_write_byteenable;                                    // nios2_dma:m_write_byteenable -> mm_interconnect_0:nios2_dma_m_write_byteenable
	wire         nios2_dma_m_write_write;                                         // nios2_dma:m_write_write -> mm_interconnect_0:nios2_dma_m_write_write
	wire  [31:0] nios2_dma_m_write_writedata;                                     // nios2_dma:m_write_writedata -> mm_interconnect_0:nios2_dma_m_write_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                           // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [27:0] nios2_cpu_instruction_master_address;                            // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                               // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_chipselect -> nios2_jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_readdata;    // nios2_jtag_uart:av_readdata -> mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_waitrequest; // nios2_jtag_uart:av_waitrequest -> mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_address -> nios2_jtag_uart:av_address
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_read -> nios2_jtag_uart:av_read_n
	wire         mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_write -> nios2_jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:nios2_jtag_uart_avalon_jtag_slave_writedata -> nios2_jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_eth1_mdio_avalon_slave_readdata;               // eth1_mdio:avalon_slave_readdata -> mm_interconnect_0:eth1_mdio_avalon_slave_readdata
	wire         mm_interconnect_0_eth1_mdio_avalon_slave_waitrequest;            // eth1_mdio:avalon_slave_waitrequest -> mm_interconnect_0:eth1_mdio_avalon_slave_waitrequest
	wire   [4:0] mm_interconnect_0_eth1_mdio_avalon_slave_address;                // mm_interconnect_0:eth1_mdio_avalon_slave_address -> eth1_mdio:avalon_slave_address
	wire         mm_interconnect_0_eth1_mdio_avalon_slave_read;                   // mm_interconnect_0:eth1_mdio_avalon_slave_read -> eth1_mdio:avalon_slave_read
	wire         mm_interconnect_0_eth1_mdio_avalon_slave_write;                  // mm_interconnect_0:eth1_mdio_avalon_slave_write -> eth1_mdio:avalon_slave_write
	wire  [31:0] mm_interconnect_0_eth1_mdio_avalon_slave_writedata;              // mm_interconnect_0:eth1_mdio_avalon_slave_writedata -> eth1_mdio:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_eth0_mdio_avalon_slave_readdata;               // eth0_mdio:avalon_slave_readdata -> mm_interconnect_0:eth0_mdio_avalon_slave_readdata
	wire         mm_interconnect_0_eth0_mdio_avalon_slave_waitrequest;            // eth0_mdio:avalon_slave_waitrequest -> mm_interconnect_0:eth0_mdio_avalon_slave_waitrequest
	wire   [4:0] mm_interconnect_0_eth0_mdio_avalon_slave_address;                // mm_interconnect_0:eth0_mdio_avalon_slave_address -> eth0_mdio:avalon_slave_address
	wire         mm_interconnect_0_eth0_mdio_avalon_slave_read;                   // mm_interconnect_0:eth0_mdio_avalon_slave_read -> eth0_mdio:avalon_slave_read
	wire         mm_interconnect_0_eth0_mdio_avalon_slave_write;                  // mm_interconnect_0:eth0_mdio_avalon_slave_write -> eth0_mdio:avalon_slave_write
	wire  [31:0] mm_interconnect_0_eth0_mdio_avalon_slave_writedata;              // mm_interconnect_0:eth0_mdio_avalon_slave_writedata -> eth0_mdio:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_sram_multiplexer_avl_readdata;                 // sram_multiplexer:AVL_READDATA -> mm_interconnect_0:sram_multiplexer_avl_readdata
	wire  [19:0] mm_interconnect_0_sram_multiplexer_avl_address;                  // mm_interconnect_0:sram_multiplexer_avl_address -> sram_multiplexer:AVL_ADDR
	wire         mm_interconnect_0_sram_multiplexer_avl_read;                     // mm_interconnect_0:sram_multiplexer_avl_read -> sram_multiplexer:AVL_READ
	wire         mm_interconnect_0_sram_multiplexer_avl_write;                    // mm_interconnect_0:sram_multiplexer_avl_write -> sram_multiplexer:AVL_WRITE
	wire  [31:0] mm_interconnect_0_sram_multiplexer_avl_writedata;                // mm_interconnect_0:sram_multiplexer_avl_writedata -> sram_multiplexer:AVL_WRITEDATA
	wire  [31:0] mm_interconnect_0_vga_sprite_params_avl_readdata;                // vga_sprite_params:AVL_READDATA -> mm_interconnect_0:vga_sprite_params_avl_readdata
	wire   [7:0] mm_interconnect_0_vga_sprite_params_avl_address;                 // mm_interconnect_0:vga_sprite_params_avl_address -> vga_sprite_params:AVL_ADDR
	wire         mm_interconnect_0_vga_sprite_params_avl_read;                    // mm_interconnect_0:vga_sprite_params_avl_read -> vga_sprite_params:AVL_READ
	wire         mm_interconnect_0_vga_sprite_params_avl_write;                   // mm_interconnect_0:vga_sprite_params_avl_write -> vga_sprite_params:AVL_WRITE
	wire  [31:0] mm_interconnect_0_vga_sprite_params_avl_writedata;               // mm_interconnect_0:vga_sprite_params_avl_writedata -> vga_sprite_params:AVL_WRITEDATA
	wire  [31:0] mm_interconnect_0_nios2_sysid_control_slave_readdata;            // nios2_sysid:readdata -> mm_interconnect_0:nios2_sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_nios2_sysid_control_slave_address;             // mm_interconnect_0:nios2_sysid_control_slave_address -> nios2_sysid:address
	wire         mm_interconnect_0_eth0_rx_dma_csr_chipselect;                    // mm_interconnect_0:eth0_rx_dma_csr_chipselect -> eth0_rx_dma:csr_chipselect
	wire  [31:0] mm_interconnect_0_eth0_rx_dma_csr_readdata;                      // eth0_rx_dma:csr_readdata -> mm_interconnect_0:eth0_rx_dma_csr_readdata
	wire   [3:0] mm_interconnect_0_eth0_rx_dma_csr_address;                       // mm_interconnect_0:eth0_rx_dma_csr_address -> eth0_rx_dma:csr_address
	wire         mm_interconnect_0_eth0_rx_dma_csr_read;                          // mm_interconnect_0:eth0_rx_dma_csr_read -> eth0_rx_dma:csr_read
	wire         mm_interconnect_0_eth0_rx_dma_csr_write;                         // mm_interconnect_0:eth0_rx_dma_csr_write -> eth0_rx_dma:csr_write
	wire  [31:0] mm_interconnect_0_eth0_rx_dma_csr_writedata;                     // mm_interconnect_0:eth0_rx_dma_csr_writedata -> eth0_rx_dma:csr_writedata
	wire         mm_interconnect_0_eth0_tx_dma_csr_chipselect;                    // mm_interconnect_0:eth0_tx_dma_csr_chipselect -> eth0_tx_dma:csr_chipselect
	wire  [31:0] mm_interconnect_0_eth0_tx_dma_csr_readdata;                      // eth0_tx_dma:csr_readdata -> mm_interconnect_0:eth0_tx_dma_csr_readdata
	wire   [3:0] mm_interconnect_0_eth0_tx_dma_csr_address;                       // mm_interconnect_0:eth0_tx_dma_csr_address -> eth0_tx_dma:csr_address
	wire         mm_interconnect_0_eth0_tx_dma_csr_read;                          // mm_interconnect_0:eth0_tx_dma_csr_read -> eth0_tx_dma:csr_read
	wire         mm_interconnect_0_eth0_tx_dma_csr_write;                         // mm_interconnect_0:eth0_tx_dma_csr_write -> eth0_tx_dma:csr_write
	wire  [31:0] mm_interconnect_0_eth0_tx_dma_csr_writedata;                     // mm_interconnect_0:eth0_tx_dma_csr_writedata -> eth0_tx_dma:csr_writedata
	wire         mm_interconnect_0_eth1_rx_dma_csr_chipselect;                    // mm_interconnect_0:eth1_rx_dma_csr_chipselect -> eth1_rx_dma:csr_chipselect
	wire  [31:0] mm_interconnect_0_eth1_rx_dma_csr_readdata;                      // eth1_rx_dma:csr_readdata -> mm_interconnect_0:eth1_rx_dma_csr_readdata
	wire   [3:0] mm_interconnect_0_eth1_rx_dma_csr_address;                       // mm_interconnect_0:eth1_rx_dma_csr_address -> eth1_rx_dma:csr_address
	wire         mm_interconnect_0_eth1_rx_dma_csr_read;                          // mm_interconnect_0:eth1_rx_dma_csr_read -> eth1_rx_dma:csr_read
	wire         mm_interconnect_0_eth1_rx_dma_csr_write;                         // mm_interconnect_0:eth1_rx_dma_csr_write -> eth1_rx_dma:csr_write
	wire  [31:0] mm_interconnect_0_eth1_rx_dma_csr_writedata;                     // mm_interconnect_0:eth1_rx_dma_csr_writedata -> eth1_rx_dma:csr_writedata
	wire         mm_interconnect_0_eth1_tx_dma_csr_chipselect;                    // mm_interconnect_0:eth1_tx_dma_csr_chipselect -> eth1_tx_dma:csr_chipselect
	wire  [31:0] mm_interconnect_0_eth1_tx_dma_csr_readdata;                      // eth1_tx_dma:csr_readdata -> mm_interconnect_0:eth1_tx_dma_csr_readdata
	wire   [3:0] mm_interconnect_0_eth1_tx_dma_csr_address;                       // mm_interconnect_0:eth1_tx_dma_csr_address -> eth1_tx_dma:csr_address
	wire         mm_interconnect_0_eth1_tx_dma_csr_read;                          // mm_interconnect_0:eth1_tx_dma_csr_read -> eth1_tx_dma:csr_read
	wire         mm_interconnect_0_eth1_tx_dma_csr_write;                         // mm_interconnect_0:eth1_tx_dma_csr_write -> eth1_tx_dma:csr_write
	wire  [31:0] mm_interconnect_0_eth1_tx_dma_csr_writedata;                     // mm_interconnect_0:eth1_tx_dma_csr_writedata -> eth1_tx_dma:csr_writedata
	wire         mm_interconnect_0_nios2_dma_csr_chipselect;                      // mm_interconnect_0:nios2_dma_csr_chipselect -> nios2_dma:csr_chipselect
	wire  [31:0] mm_interconnect_0_nios2_dma_csr_readdata;                        // nios2_dma:csr_readdata -> mm_interconnect_0:nios2_dma_csr_readdata
	wire   [3:0] mm_interconnect_0_nios2_dma_csr_address;                         // mm_interconnect_0:nios2_dma_csr_address -> nios2_dma:csr_address
	wire         mm_interconnect_0_nios2_dma_csr_read;                            // mm_interconnect_0:nios2_dma_csr_read -> nios2_dma:csr_read
	wire         mm_interconnect_0_nios2_dma_csr_write;                           // mm_interconnect_0:nios2_dma_csr_write -> nios2_dma:csr_write
	wire  [31:0] mm_interconnect_0_nios2_dma_csr_writedata;                       // mm_interconnect_0:nios2_dma_csr_writedata -> nios2_dma:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;            // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;         // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;             // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;                // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;               // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_nios2_pll_pll_slave_readdata;                  // nios2_pll:readdata -> mm_interconnect_0:nios2_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_nios2_pll_pll_slave_address;                   // mm_interconnect_0:nios2_pll_pll_slave_address -> nios2_pll:address
	wire         mm_interconnect_0_nios2_pll_pll_slave_read;                      // mm_interconnect_0:nios2_pll_pll_slave_read -> nios2_pll:read
	wire         mm_interconnect_0_nios2_pll_pll_slave_write;                     // mm_interconnect_0:nios2_pll_pll_slave_write -> nios2_pll:write
	wire  [31:0] mm_interconnect_0_nios2_pll_pll_slave_writedata;                 // mm_interconnect_0:nios2_pll_pll_slave_writedata -> nios2_pll:writedata
	wire         mm_interconnect_0_nios2_onchip_mem_s1_chipselect;                // mm_interconnect_0:nios2_onchip_mem_s1_chipselect -> nios2_onchip_mem:chipselect
	wire  [31:0] mm_interconnect_0_nios2_onchip_mem_s1_readdata;                  // nios2_onchip_mem:readdata -> mm_interconnect_0:nios2_onchip_mem_s1_readdata
	wire  [15:0] mm_interconnect_0_nios2_onchip_mem_s1_address;                   // mm_interconnect_0:nios2_onchip_mem_s1_address -> nios2_onchip_mem:address
	wire   [3:0] mm_interconnect_0_nios2_onchip_mem_s1_byteenable;                // mm_interconnect_0:nios2_onchip_mem_s1_byteenable -> nios2_onchip_mem:byteenable
	wire         mm_interconnect_0_nios2_onchip_mem_s1_write;                     // mm_interconnect_0:nios2_onchip_mem_s1_write -> nios2_onchip_mem:write
	wire  [31:0] mm_interconnect_0_nios2_onchip_mem_s1_writedata;                 // mm_interconnect_0:nios2_onchip_mem_s1_writedata -> nios2_onchip_mem:writedata
	wire         mm_interconnect_0_nios2_onchip_mem_s1_clken;                     // mm_interconnect_0:nios2_onchip_mem_s1_clken -> nios2_onchip_mem:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                           // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                             // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                          // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                              // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                 // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                           // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                        // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                            // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_io_led_red_s1_chipselect;                      // mm_interconnect_0:io_led_red_s1_chipselect -> io_led_red:chipselect
	wire  [31:0] mm_interconnect_0_io_led_red_s1_readdata;                        // io_led_red:readdata -> mm_interconnect_0:io_led_red_s1_readdata
	wire   [2:0] mm_interconnect_0_io_led_red_s1_address;                         // mm_interconnect_0:io_led_red_s1_address -> io_led_red:address
	wire         mm_interconnect_0_io_led_red_s1_write;                           // mm_interconnect_0:io_led_red_s1_write -> io_led_red:write_n
	wire  [31:0] mm_interconnect_0_io_led_red_s1_writedata;                       // mm_interconnect_0:io_led_red_s1_writedata -> io_led_red:writedata
	wire         mm_interconnect_0_nios2_timer_s1_chipselect;                     // mm_interconnect_0:nios2_timer_s1_chipselect -> nios2_timer:chipselect
	wire  [15:0] mm_interconnect_0_nios2_timer_s1_readdata;                       // nios2_timer:readdata -> mm_interconnect_0:nios2_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_nios2_timer_s1_address;                        // mm_interconnect_0:nios2_timer_s1_address -> nios2_timer:address
	wire         mm_interconnect_0_nios2_timer_s1_write;                          // mm_interconnect_0:nios2_timer_s1_write -> nios2_timer:write_n
	wire  [15:0] mm_interconnect_0_nios2_timer_s1_writedata;                      // mm_interconnect_0:nios2_timer_s1_writedata -> nios2_timer:writedata
	wire  [31:0] mm_interconnect_0_io_keys_s1_readdata;                           // io_keys:readdata -> mm_interconnect_0:io_keys_s1_readdata
	wire   [1:0] mm_interconnect_0_io_keys_s1_address;                            // mm_interconnect_0:io_keys_s1_address -> io_keys:address
	wire  [31:0] mm_interconnect_0_io_switches_s1_readdata;                       // io_switches:readdata -> mm_interconnect_0:io_switches_s1_readdata
	wire   [1:0] mm_interconnect_0_io_switches_s1_address;                        // mm_interconnect_0:io_switches_s1_address -> io_switches:address
	wire         mm_interconnect_0_io_led_green_s1_chipselect;                    // mm_interconnect_0:io_led_green_s1_chipselect -> io_led_green:chipselect
	wire  [31:0] mm_interconnect_0_io_led_green_s1_readdata;                      // io_led_green:readdata -> mm_interconnect_0:io_led_green_s1_readdata
	wire   [2:0] mm_interconnect_0_io_led_green_s1_address;                       // mm_interconnect_0:io_led_green_s1_address -> io_led_green:address
	wire         mm_interconnect_0_io_led_green_s1_write;                         // mm_interconnect_0:io_led_green_s1_write -> io_led_green:write_n
	wire  [31:0] mm_interconnect_0_io_led_green_s1_writedata;                     // mm_interconnect_0:io_led_green_s1_writedata -> io_led_green:writedata
	wire         mm_interconnect_0_io_hex_s1_chipselect;                          // mm_interconnect_0:io_hex_s1_chipselect -> io_hex:chipselect
	wire  [31:0] mm_interconnect_0_io_hex_s1_readdata;                            // io_hex:readdata -> mm_interconnect_0:io_hex_s1_readdata
	wire   [2:0] mm_interconnect_0_io_hex_s1_address;                             // mm_interconnect_0:io_hex_s1_address -> io_hex:address
	wire         mm_interconnect_0_io_hex_s1_write;                               // mm_interconnect_0:io_hex_s1_write -> io_hex:write_n
	wire  [31:0] mm_interconnect_0_io_hex_s1_writedata;                           // mm_interconnect_0:io_hex_s1_writedata -> io_hex:writedata
	wire         mm_interconnect_0_vga_sprite_0_s1_chipselect;                    // mm_interconnect_0:vga_sprite_0_s1_chipselect -> vga_sprite_0:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_0_s1_readdata;                      // vga_sprite_0:readdata -> mm_interconnect_0:vga_sprite_0_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_0_s1_address;                       // mm_interconnect_0:vga_sprite_0_s1_address -> vga_sprite_0:address
	wire   [3:0] mm_interconnect_0_vga_sprite_0_s1_byteenable;                    // mm_interconnect_0:vga_sprite_0_s1_byteenable -> vga_sprite_0:byteenable
	wire         mm_interconnect_0_vga_sprite_0_s1_write;                         // mm_interconnect_0:vga_sprite_0_s1_write -> vga_sprite_0:write
	wire  [31:0] mm_interconnect_0_vga_sprite_0_s1_writedata;                     // mm_interconnect_0:vga_sprite_0_s1_writedata -> vga_sprite_0:writedata
	wire         mm_interconnect_0_vga_sprite_0_s1_clken;                         // mm_interconnect_0:vga_sprite_0_s1_clken -> vga_sprite_0:clken
	wire         mm_interconnect_0_vga_sprite_1_s1_chipselect;                    // mm_interconnect_0:vga_sprite_1_s1_chipselect -> vga_sprite_1:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_1_s1_readdata;                      // vga_sprite_1:readdata -> mm_interconnect_0:vga_sprite_1_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_1_s1_address;                       // mm_interconnect_0:vga_sprite_1_s1_address -> vga_sprite_1:address
	wire   [3:0] mm_interconnect_0_vga_sprite_1_s1_byteenable;                    // mm_interconnect_0:vga_sprite_1_s1_byteenable -> vga_sprite_1:byteenable
	wire         mm_interconnect_0_vga_sprite_1_s1_write;                         // mm_interconnect_0:vga_sprite_1_s1_write -> vga_sprite_1:write
	wire  [31:0] mm_interconnect_0_vga_sprite_1_s1_writedata;                     // mm_interconnect_0:vga_sprite_1_s1_writedata -> vga_sprite_1:writedata
	wire         mm_interconnect_0_vga_sprite_1_s1_clken;                         // mm_interconnect_0:vga_sprite_1_s1_clken -> vga_sprite_1:clken
	wire         mm_interconnect_0_vga_sprite_2_s1_chipselect;                    // mm_interconnect_0:vga_sprite_2_s1_chipselect -> vga_sprite_2:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_2_s1_readdata;                      // vga_sprite_2:readdata -> mm_interconnect_0:vga_sprite_2_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_2_s1_address;                       // mm_interconnect_0:vga_sprite_2_s1_address -> vga_sprite_2:address
	wire   [3:0] mm_interconnect_0_vga_sprite_2_s1_byteenable;                    // mm_interconnect_0:vga_sprite_2_s1_byteenable -> vga_sprite_2:byteenable
	wire         mm_interconnect_0_vga_sprite_2_s1_write;                         // mm_interconnect_0:vga_sprite_2_s1_write -> vga_sprite_2:write
	wire  [31:0] mm_interconnect_0_vga_sprite_2_s1_writedata;                     // mm_interconnect_0:vga_sprite_2_s1_writedata -> vga_sprite_2:writedata
	wire         mm_interconnect_0_vga_sprite_2_s1_clken;                         // mm_interconnect_0:vga_sprite_2_s1_clken -> vga_sprite_2:clken
	wire         mm_interconnect_0_vga_sprite_3_s1_chipselect;                    // mm_interconnect_0:vga_sprite_3_s1_chipselect -> vga_sprite_3:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_3_s1_readdata;                      // vga_sprite_3:readdata -> mm_interconnect_0:vga_sprite_3_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_3_s1_address;                       // mm_interconnect_0:vga_sprite_3_s1_address -> vga_sprite_3:address
	wire   [3:0] mm_interconnect_0_vga_sprite_3_s1_byteenable;                    // mm_interconnect_0:vga_sprite_3_s1_byteenable -> vga_sprite_3:byteenable
	wire         mm_interconnect_0_vga_sprite_3_s1_write;                         // mm_interconnect_0:vga_sprite_3_s1_write -> vga_sprite_3:write
	wire  [31:0] mm_interconnect_0_vga_sprite_3_s1_writedata;                     // mm_interconnect_0:vga_sprite_3_s1_writedata -> vga_sprite_3:writedata
	wire         mm_interconnect_0_vga_sprite_3_s1_clken;                         // mm_interconnect_0:vga_sprite_3_s1_clken -> vga_sprite_3:clken
	wire  [31:0] mm_interconnect_0_io_vga_sync_s1_readdata;                       // io_vga_sync:readdata -> mm_interconnect_0:io_vga_sync_s1_readdata
	wire   [1:0] mm_interconnect_0_io_vga_sync_s1_address;                        // mm_interconnect_0:io_vga_sync_s1_address -> io_vga_sync:address
	wire         mm_interconnect_0_vga_sprite_4_s1_chipselect;                    // mm_interconnect_0:vga_sprite_4_s1_chipselect -> vga_sprite_4:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_4_s1_readdata;                      // vga_sprite_4:readdata -> mm_interconnect_0:vga_sprite_4_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_4_s1_address;                       // mm_interconnect_0:vga_sprite_4_s1_address -> vga_sprite_4:address
	wire   [3:0] mm_interconnect_0_vga_sprite_4_s1_byteenable;                    // mm_interconnect_0:vga_sprite_4_s1_byteenable -> vga_sprite_4:byteenable
	wire         mm_interconnect_0_vga_sprite_4_s1_write;                         // mm_interconnect_0:vga_sprite_4_s1_write -> vga_sprite_4:write
	wire  [31:0] mm_interconnect_0_vga_sprite_4_s1_writedata;                     // mm_interconnect_0:vga_sprite_4_s1_writedata -> vga_sprite_4:writedata
	wire         mm_interconnect_0_vga_sprite_4_s1_clken;                         // mm_interconnect_0:vga_sprite_4_s1_clken -> vga_sprite_4:clken
	wire         mm_interconnect_0_vga_sprite_5_s1_chipselect;                    // mm_interconnect_0:vga_sprite_5_s1_chipselect -> vga_sprite_5:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_5_s1_readdata;                      // vga_sprite_5:readdata -> mm_interconnect_0:vga_sprite_5_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_5_s1_address;                       // mm_interconnect_0:vga_sprite_5_s1_address -> vga_sprite_5:address
	wire   [3:0] mm_interconnect_0_vga_sprite_5_s1_byteenable;                    // mm_interconnect_0:vga_sprite_5_s1_byteenable -> vga_sprite_5:byteenable
	wire         mm_interconnect_0_vga_sprite_5_s1_write;                         // mm_interconnect_0:vga_sprite_5_s1_write -> vga_sprite_5:write
	wire  [31:0] mm_interconnect_0_vga_sprite_5_s1_writedata;                     // mm_interconnect_0:vga_sprite_5_s1_writedata -> vga_sprite_5:writedata
	wire         mm_interconnect_0_vga_sprite_5_s1_clken;                         // mm_interconnect_0:vga_sprite_5_s1_clken -> vga_sprite_5:clken
	wire         mm_interconnect_0_vga_sprite_6_s1_chipselect;                    // mm_interconnect_0:vga_sprite_6_s1_chipselect -> vga_sprite_6:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_6_s1_readdata;                      // vga_sprite_6:readdata -> mm_interconnect_0:vga_sprite_6_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_6_s1_address;                       // mm_interconnect_0:vga_sprite_6_s1_address -> vga_sprite_6:address
	wire   [3:0] mm_interconnect_0_vga_sprite_6_s1_byteenable;                    // mm_interconnect_0:vga_sprite_6_s1_byteenable -> vga_sprite_6:byteenable
	wire         mm_interconnect_0_vga_sprite_6_s1_write;                         // mm_interconnect_0:vga_sprite_6_s1_write -> vga_sprite_6:write
	wire  [31:0] mm_interconnect_0_vga_sprite_6_s1_writedata;                     // mm_interconnect_0:vga_sprite_6_s1_writedata -> vga_sprite_6:writedata
	wire         mm_interconnect_0_vga_sprite_6_s1_clken;                         // mm_interconnect_0:vga_sprite_6_s1_clken -> vga_sprite_6:clken
	wire         mm_interconnect_0_vga_sprite_7_s1_chipselect;                    // mm_interconnect_0:vga_sprite_7_s1_chipselect -> vga_sprite_7:chipselect
	wire  [31:0] mm_interconnect_0_vga_sprite_7_s1_readdata;                      // vga_sprite_7:readdata -> mm_interconnect_0:vga_sprite_7_s1_readdata
	wire   [9:0] mm_interconnect_0_vga_sprite_7_s1_address;                       // mm_interconnect_0:vga_sprite_7_s1_address -> vga_sprite_7:address
	wire   [3:0] mm_interconnect_0_vga_sprite_7_s1_byteenable;                    // mm_interconnect_0:vga_sprite_7_s1_byteenable -> vga_sprite_7:byteenable
	wire         mm_interconnect_0_vga_sprite_7_s1_write;                         // mm_interconnect_0:vga_sprite_7_s1_write -> vga_sprite_7:write
	wire  [31:0] mm_interconnect_0_vga_sprite_7_s1_writedata;                     // mm_interconnect_0:vga_sprite_7_s1_writedata -> vga_sprite_7:writedata
	wire         mm_interconnect_0_vga_sprite_7_s1_clken;                         // mm_interconnect_0:vga_sprite_7_s1_clken -> vga_sprite_7:clken
	wire         mm_interconnect_0_audio_mem_s1_chipselect;                       // mm_interconnect_0:audio_mem_s1_chipselect -> audio_mem:chipselect
	wire  [31:0] mm_interconnect_0_audio_mem_s1_readdata;                         // audio_mem:readdata -> mm_interconnect_0:audio_mem_s1_readdata
	wire  [11:0] mm_interconnect_0_audio_mem_s1_address;                          // mm_interconnect_0:audio_mem_s1_address -> audio_mem:address
	wire   [3:0] mm_interconnect_0_audio_mem_s1_byteenable;                       // mm_interconnect_0:audio_mem_s1_byteenable -> audio_mem:byteenable
	wire         mm_interconnect_0_audio_mem_s1_write;                            // mm_interconnect_0:audio_mem_s1_write -> audio_mem:write
	wire  [31:0] mm_interconnect_0_audio_mem_s1_writedata;                        // mm_interconnect_0:audio_mem_s1_writedata -> audio_mem:writedata
	wire         mm_interconnect_0_audio_mem_s1_clken;                            // mm_interconnect_0:audio_mem_s1_clken -> audio_mem:clken
	wire         mm_interconnect_0_audio_position_end_s1_chipselect;              // mm_interconnect_0:audio_position_end_s1_chipselect -> audio_position_end:chipselect
	wire  [31:0] mm_interconnect_0_audio_position_end_s1_readdata;                // audio_position_end:readdata -> mm_interconnect_0:audio_position_end_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_position_end_s1_address;                 // mm_interconnect_0:audio_position_end_s1_address -> audio_position_end:address
	wire         mm_interconnect_0_audio_position_end_s1_write;                   // mm_interconnect_0:audio_position_end_s1_write -> audio_position_end:write_n
	wire  [31:0] mm_interconnect_0_audio_position_end_s1_writedata;               // mm_interconnect_0:audio_position_end_s1_writedata -> audio_position_end:writedata
	wire  [31:0] mm_interconnect_0_audio_position_s1_readdata;                    // audio_position:readdata -> mm_interconnect_0:audio_position_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_position_s1_address;                     // mm_interconnect_0:audio_position_s1_address -> audio_position:address
	wire         mm_interconnect_0_vga_background_offset_s1_chipselect;           // mm_interconnect_0:vga_background_offset_s1_chipselect -> vga_background_offset:chipselect
	wire  [31:0] mm_interconnect_0_vga_background_offset_s1_readdata;             // vga_background_offset:readdata -> mm_interconnect_0:vga_background_offset_s1_readdata
	wire   [1:0] mm_interconnect_0_vga_background_offset_s1_address;              // mm_interconnect_0:vga_background_offset_s1_address -> vga_background_offset:address
	wire         mm_interconnect_0_vga_background_offset_s1_write;                // mm_interconnect_0:vga_background_offset_s1_write -> vga_background_offset:write_n
	wire  [31:0] mm_interconnect_0_vga_background_offset_s1_writedata;            // mm_interconnect_0:vga_background_offset_s1_writedata -> vga_background_offset:writedata
	wire         mm_interconnect_0_usb_keycode_s2_chipselect;                     // mm_interconnect_0:usb_keycode_s2_chipselect -> usb_keycode:chipselect2
	wire  [31:0] mm_interconnect_0_usb_keycode_s2_readdata;                       // usb_keycode:readdata2 -> mm_interconnect_0:usb_keycode_s2_readdata
	wire   [7:0] mm_interconnect_0_usb_keycode_s2_address;                        // mm_interconnect_0:usb_keycode_s2_address -> usb_keycode:address2
	wire   [3:0] mm_interconnect_0_usb_keycode_s2_byteenable;                     // mm_interconnect_0:usb_keycode_s2_byteenable -> usb_keycode:byteenable2
	wire         mm_interconnect_0_usb_keycode_s2_write;                          // mm_interconnect_0:usb_keycode_s2_write -> usb_keycode:write2
	wire  [31:0] mm_interconnect_0_usb_keycode_s2_writedata;                      // mm_interconnect_0:usb_keycode_s2_writedata -> usb_keycode:writedata2
	wire         mm_interconnect_0_usb_keycode_s2_clken;                          // mm_interconnect_0:usb_keycode_s2_clken -> usb_keycode:clken2
	wire  [31:0] usb_nios2_cpu_data_master_readdata;                              // mm_interconnect_1:usb_nios2_cpu_data_master_readdata -> usb_nios2_cpu:d_readdata
	wire         usb_nios2_cpu_data_master_waitrequest;                           // mm_interconnect_1:usb_nios2_cpu_data_master_waitrequest -> usb_nios2_cpu:d_waitrequest
	wire         usb_nios2_cpu_data_master_debugaccess;                           // usb_nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:usb_nios2_cpu_data_master_debugaccess
	wire  [16:0] usb_nios2_cpu_data_master_address;                               // usb_nios2_cpu:d_address -> mm_interconnect_1:usb_nios2_cpu_data_master_address
	wire   [3:0] usb_nios2_cpu_data_master_byteenable;                            // usb_nios2_cpu:d_byteenable -> mm_interconnect_1:usb_nios2_cpu_data_master_byteenable
	wire         usb_nios2_cpu_data_master_read;                                  // usb_nios2_cpu:d_read -> mm_interconnect_1:usb_nios2_cpu_data_master_read
	wire         usb_nios2_cpu_data_master_write;                                 // usb_nios2_cpu:d_write -> mm_interconnect_1:usb_nios2_cpu_data_master_write
	wire  [31:0] usb_nios2_cpu_data_master_writedata;                             // usb_nios2_cpu:d_writedata -> mm_interconnect_1:usb_nios2_cpu_data_master_writedata
	wire  [31:0] usb_nios2_cpu_instruction_master_readdata;                       // mm_interconnect_1:usb_nios2_cpu_instruction_master_readdata -> usb_nios2_cpu:i_readdata
	wire         usb_nios2_cpu_instruction_master_waitrequest;                    // mm_interconnect_1:usb_nios2_cpu_instruction_master_waitrequest -> usb_nios2_cpu:i_waitrequest
	wire  [16:0] usb_nios2_cpu_instruction_master_address;                        // usb_nios2_cpu:i_address -> mm_interconnect_1:usb_nios2_cpu_instruction_master_address
	wire         usb_nios2_cpu_instruction_master_read;                           // usb_nios2_cpu:i_read -> mm_interconnect_1:usb_nios2_cpu_instruction_master_read
	wire         mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_1:usb_jtag_uart_avalon_jtag_slave_chipselect -> usb_jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_readdata;      // usb_jtag_uart:av_readdata -> mm_interconnect_1:usb_jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_waitrequest;   // usb_jtag_uart:av_waitrequest -> mm_interconnect_1:usb_jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_address;       // mm_interconnect_1:usb_jtag_uart_avalon_jtag_slave_address -> usb_jtag_uart:av_address
	wire         mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_read;          // mm_interconnect_1:usb_jtag_uart_avalon_jtag_slave_read -> usb_jtag_uart:av_read_n
	wire         mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_write;         // mm_interconnect_1:usb_jtag_uart_avalon_jtag_slave_write -> usb_jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_writedata;     // mm_interconnect_1:usb_jtag_uart_avalon_jtag_slave_writedata -> usb_jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_usb_nios2_sysid_control_slave_readdata;        // usb_nios2_sysid:readdata -> mm_interconnect_1:usb_nios2_sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_usb_nios2_sysid_control_slave_address;         // mm_interconnect_1:usb_nios2_sysid_control_slave_address -> usb_nios2_sysid:address
	wire  [31:0] mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_readdata;        // usb_nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_waitrequest;     // usb_nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_debugaccess;     // mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_debugaccess -> usb_nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_address;         // mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_address -> usb_nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_read;            // mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_read -> usb_nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_byteenable;      // mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_byteenable -> usb_nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_write;           // mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_write -> usb_nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_writedata;       // mm_interconnect_1:usb_nios2_cpu_debug_mem_slave_writedata -> usb_nios2_cpu:debug_mem_slave_writedata
	wire         mm_interconnect_1_usb_nios2_onchip_mem_s1_chipselect;            // mm_interconnect_1:usb_nios2_onchip_mem_s1_chipselect -> usb_nios2_onchip_mem:chipselect
	wire  [31:0] mm_interconnect_1_usb_nios2_onchip_mem_s1_readdata;              // usb_nios2_onchip_mem:readdata -> mm_interconnect_1:usb_nios2_onchip_mem_s1_readdata
	wire  [11:0] mm_interconnect_1_usb_nios2_onchip_mem_s1_address;               // mm_interconnect_1:usb_nios2_onchip_mem_s1_address -> usb_nios2_onchip_mem:address
	wire   [3:0] mm_interconnect_1_usb_nios2_onchip_mem_s1_byteenable;            // mm_interconnect_1:usb_nios2_onchip_mem_s1_byteenable -> usb_nios2_onchip_mem:byteenable
	wire         mm_interconnect_1_usb_nios2_onchip_mem_s1_write;                 // mm_interconnect_1:usb_nios2_onchip_mem_s1_write -> usb_nios2_onchip_mem:write
	wire  [31:0] mm_interconnect_1_usb_nios2_onchip_mem_s1_writedata;             // mm_interconnect_1:usb_nios2_onchip_mem_s1_writedata -> usb_nios2_onchip_mem:writedata
	wire         mm_interconnect_1_usb_nios2_onchip_mem_s1_clken;                 // mm_interconnect_1:usb_nios2_onchip_mem_s1_clken -> usb_nios2_onchip_mem:clken
	wire         mm_interconnect_1_usb_hpi_reset_s1_chipselect;                   // mm_interconnect_1:usb_hpi_reset_s1_chipselect -> usb_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_1_usb_hpi_reset_s1_readdata;                     // usb_hpi_reset:readdata -> mm_interconnect_1:usb_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_1_usb_hpi_reset_s1_address;                      // mm_interconnect_1:usb_hpi_reset_s1_address -> usb_hpi_reset:address
	wire         mm_interconnect_1_usb_hpi_reset_s1_write;                        // mm_interconnect_1:usb_hpi_reset_s1_write -> usb_hpi_reset:write_n
	wire  [31:0] mm_interconnect_1_usb_hpi_reset_s1_writedata;                    // mm_interconnect_1:usb_hpi_reset_s1_writedata -> usb_hpi_reset:writedata
	wire         mm_interconnect_1_usb_hpi_cs_s1_chipselect;                      // mm_interconnect_1:usb_hpi_cs_s1_chipselect -> usb_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_1_usb_hpi_cs_s1_readdata;                        // usb_hpi_cs:readdata -> mm_interconnect_1:usb_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_1_usb_hpi_cs_s1_address;                         // mm_interconnect_1:usb_hpi_cs_s1_address -> usb_hpi_cs:address
	wire         mm_interconnect_1_usb_hpi_cs_s1_write;                           // mm_interconnect_1:usb_hpi_cs_s1_write -> usb_hpi_cs:write_n
	wire  [31:0] mm_interconnect_1_usb_hpi_cs_s1_writedata;                       // mm_interconnect_1:usb_hpi_cs_s1_writedata -> usb_hpi_cs:writedata
	wire         mm_interconnect_1_usb_hpi_w_s1_chipselect;                       // mm_interconnect_1:usb_hpi_w_s1_chipselect -> usb_hpi_w:chipselect
	wire  [31:0] mm_interconnect_1_usb_hpi_w_s1_readdata;                         // usb_hpi_w:readdata -> mm_interconnect_1:usb_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_1_usb_hpi_w_s1_address;                          // mm_interconnect_1:usb_hpi_w_s1_address -> usb_hpi_w:address
	wire         mm_interconnect_1_usb_hpi_w_s1_write;                            // mm_interconnect_1:usb_hpi_w_s1_write -> usb_hpi_w:write_n
	wire  [31:0] mm_interconnect_1_usb_hpi_w_s1_writedata;                        // mm_interconnect_1:usb_hpi_w_s1_writedata -> usb_hpi_w:writedata
	wire         mm_interconnect_1_usb_hpi_r_s1_chipselect;                       // mm_interconnect_1:usb_hpi_r_s1_chipselect -> usb_hpi_r:chipselect
	wire  [31:0] mm_interconnect_1_usb_hpi_r_s1_readdata;                         // usb_hpi_r:readdata -> mm_interconnect_1:usb_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_1_usb_hpi_r_s1_address;                          // mm_interconnect_1:usb_hpi_r_s1_address -> usb_hpi_r:address
	wire         mm_interconnect_1_usb_hpi_r_s1_write;                            // mm_interconnect_1:usb_hpi_r_s1_write -> usb_hpi_r:write_n
	wire  [31:0] mm_interconnect_1_usb_hpi_r_s1_writedata;                        // mm_interconnect_1:usb_hpi_r_s1_writedata -> usb_hpi_r:writedata
	wire         mm_interconnect_1_usb_hpi_data_s1_chipselect;                    // mm_interconnect_1:usb_hpi_data_s1_chipselect -> usb_hpi_data:chipselect
	wire  [31:0] mm_interconnect_1_usb_hpi_data_s1_readdata;                      // usb_hpi_data:readdata -> mm_interconnect_1:usb_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_1_usb_hpi_data_s1_address;                       // mm_interconnect_1:usb_hpi_data_s1_address -> usb_hpi_data:address
	wire         mm_interconnect_1_usb_hpi_data_s1_write;                         // mm_interconnect_1:usb_hpi_data_s1_write -> usb_hpi_data:write_n
	wire  [31:0] mm_interconnect_1_usb_hpi_data_s1_writedata;                     // mm_interconnect_1:usb_hpi_data_s1_writedata -> usb_hpi_data:writedata
	wire         mm_interconnect_1_usb_hpi_address_s1_chipselect;                 // mm_interconnect_1:usb_hpi_address_s1_chipselect -> usb_hpi_address:chipselect
	wire  [31:0] mm_interconnect_1_usb_hpi_address_s1_readdata;                   // usb_hpi_address:readdata -> mm_interconnect_1:usb_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_1_usb_hpi_address_s1_address;                    // mm_interconnect_1:usb_hpi_address_s1_address -> usb_hpi_address:address
	wire         mm_interconnect_1_usb_hpi_address_s1_write;                      // mm_interconnect_1:usb_hpi_address_s1_write -> usb_hpi_address:write_n
	wire  [31:0] mm_interconnect_1_usb_hpi_address_s1_writedata;                  // mm_interconnect_1:usb_hpi_address_s1_writedata -> usb_hpi_address:writedata
	wire         mm_interconnect_1_usb_keycode_s1_chipselect;                     // mm_interconnect_1:usb_keycode_s1_chipselect -> usb_keycode:chipselect
	wire  [31:0] mm_interconnect_1_usb_keycode_s1_readdata;                       // usb_keycode:readdata -> mm_interconnect_1:usb_keycode_s1_readdata
	wire   [7:0] mm_interconnect_1_usb_keycode_s1_address;                        // mm_interconnect_1:usb_keycode_s1_address -> usb_keycode:address
	wire   [3:0] mm_interconnect_1_usb_keycode_s1_byteenable;                     // mm_interconnect_1:usb_keycode_s1_byteenable -> usb_keycode:byteenable
	wire         mm_interconnect_1_usb_keycode_s1_write;                          // mm_interconnect_1:usb_keycode_s1_write -> usb_keycode:write
	wire  [31:0] mm_interconnect_1_usb_keycode_s1_writedata;                      // mm_interconnect_1:usb_keycode_s1_writedata -> usb_keycode:writedata
	wire         mm_interconnect_1_usb_keycode_s1_clken;                          // mm_interconnect_1:usb_keycode_s1_clken -> usb_keycode:clken
	wire  [31:0] eth0_rx_dma_descriptor_read_readdata;                            // mm_interconnect_2:eth0_rx_dma_descriptor_read_readdata -> eth0_rx_dma:descriptor_read_readdata
	wire         eth0_rx_dma_descriptor_read_waitrequest;                         // mm_interconnect_2:eth0_rx_dma_descriptor_read_waitrequest -> eth0_rx_dma:descriptor_read_waitrequest
	wire  [31:0] eth0_rx_dma_descriptor_read_address;                             // eth0_rx_dma:descriptor_read_address -> mm_interconnect_2:eth0_rx_dma_descriptor_read_address
	wire         eth0_rx_dma_descriptor_read_read;                                // eth0_rx_dma:descriptor_read_read -> mm_interconnect_2:eth0_rx_dma_descriptor_read_read
	wire         eth0_rx_dma_descriptor_read_readdatavalid;                       // mm_interconnect_2:eth0_rx_dma_descriptor_read_readdatavalid -> eth0_rx_dma:descriptor_read_readdatavalid
	wire  [31:0] eth0_tx_dma_descriptor_read_readdata;                            // mm_interconnect_2:eth0_tx_dma_descriptor_read_readdata -> eth0_tx_dma:descriptor_read_readdata
	wire         eth0_tx_dma_descriptor_read_waitrequest;                         // mm_interconnect_2:eth0_tx_dma_descriptor_read_waitrequest -> eth0_tx_dma:descriptor_read_waitrequest
	wire  [31:0] eth0_tx_dma_descriptor_read_address;                             // eth0_tx_dma:descriptor_read_address -> mm_interconnect_2:eth0_tx_dma_descriptor_read_address
	wire         eth0_tx_dma_descriptor_read_read;                                // eth0_tx_dma:descriptor_read_read -> mm_interconnect_2:eth0_tx_dma_descriptor_read_read
	wire         eth0_tx_dma_descriptor_read_readdatavalid;                       // mm_interconnect_2:eth0_tx_dma_descriptor_read_readdatavalid -> eth0_tx_dma:descriptor_read_readdatavalid
	wire  [31:0] eth1_rx_dma_descriptor_read_readdata;                            // mm_interconnect_2:eth1_rx_dma_descriptor_read_readdata -> eth1_rx_dma:descriptor_read_readdata
	wire         eth1_rx_dma_descriptor_read_waitrequest;                         // mm_interconnect_2:eth1_rx_dma_descriptor_read_waitrequest -> eth1_rx_dma:descriptor_read_waitrequest
	wire  [31:0] eth1_rx_dma_descriptor_read_address;                             // eth1_rx_dma:descriptor_read_address -> mm_interconnect_2:eth1_rx_dma_descriptor_read_address
	wire         eth1_rx_dma_descriptor_read_read;                                // eth1_rx_dma:descriptor_read_read -> mm_interconnect_2:eth1_rx_dma_descriptor_read_read
	wire         eth1_rx_dma_descriptor_read_readdatavalid;                       // mm_interconnect_2:eth1_rx_dma_descriptor_read_readdatavalid -> eth1_rx_dma:descriptor_read_readdatavalid
	wire  [31:0] eth1_tx_dma_descriptor_read_readdata;                            // mm_interconnect_2:eth1_tx_dma_descriptor_read_readdata -> eth1_tx_dma:descriptor_read_readdata
	wire         eth1_tx_dma_descriptor_read_waitrequest;                         // mm_interconnect_2:eth1_tx_dma_descriptor_read_waitrequest -> eth1_tx_dma:descriptor_read_waitrequest
	wire  [31:0] eth1_tx_dma_descriptor_read_address;                             // eth1_tx_dma:descriptor_read_address -> mm_interconnect_2:eth1_tx_dma_descriptor_read_address
	wire         eth1_tx_dma_descriptor_read_read;                                // eth1_tx_dma:descriptor_read_read -> mm_interconnect_2:eth1_tx_dma_descriptor_read_read
	wire         eth1_tx_dma_descriptor_read_readdatavalid;                       // mm_interconnect_2:eth1_tx_dma_descriptor_read_readdatavalid -> eth1_tx_dma:descriptor_read_readdatavalid
	wire  [31:0] nios2_dma_descriptor_read_readdata;                              // mm_interconnect_2:nios2_dma_descriptor_read_readdata -> nios2_dma:descriptor_read_readdata
	wire         nios2_dma_descriptor_read_waitrequest;                           // mm_interconnect_2:nios2_dma_descriptor_read_waitrequest -> nios2_dma:descriptor_read_waitrequest
	wire  [31:0] nios2_dma_descriptor_read_address;                               // nios2_dma:descriptor_read_address -> mm_interconnect_2:nios2_dma_descriptor_read_address
	wire         nios2_dma_descriptor_read_read;                                  // nios2_dma:descriptor_read_read -> mm_interconnect_2:nios2_dma_descriptor_read_read
	wire         nios2_dma_descriptor_read_readdatavalid;                         // mm_interconnect_2:nios2_dma_descriptor_read_readdatavalid -> nios2_dma:descriptor_read_readdatavalid
	wire         eth0_rx_dma_descriptor_write_waitrequest;                        // mm_interconnect_2:eth0_rx_dma_descriptor_write_waitrequest -> eth0_rx_dma:descriptor_write_waitrequest
	wire  [31:0] eth0_rx_dma_descriptor_write_address;                            // eth0_rx_dma:descriptor_write_address -> mm_interconnect_2:eth0_rx_dma_descriptor_write_address
	wire         eth0_rx_dma_descriptor_write_write;                              // eth0_rx_dma:descriptor_write_write -> mm_interconnect_2:eth0_rx_dma_descriptor_write_write
	wire  [31:0] eth0_rx_dma_descriptor_write_writedata;                          // eth0_rx_dma:descriptor_write_writedata -> mm_interconnect_2:eth0_rx_dma_descriptor_write_writedata
	wire         eth0_tx_dma_descriptor_write_waitrequest;                        // mm_interconnect_2:eth0_tx_dma_descriptor_write_waitrequest -> eth0_tx_dma:descriptor_write_waitrequest
	wire  [31:0] eth0_tx_dma_descriptor_write_address;                            // eth0_tx_dma:descriptor_write_address -> mm_interconnect_2:eth0_tx_dma_descriptor_write_address
	wire         eth0_tx_dma_descriptor_write_write;                              // eth0_tx_dma:descriptor_write_write -> mm_interconnect_2:eth0_tx_dma_descriptor_write_write
	wire  [31:0] eth0_tx_dma_descriptor_write_writedata;                          // eth0_tx_dma:descriptor_write_writedata -> mm_interconnect_2:eth0_tx_dma_descriptor_write_writedata
	wire         eth1_rx_dma_descriptor_write_waitrequest;                        // mm_interconnect_2:eth1_rx_dma_descriptor_write_waitrequest -> eth1_rx_dma:descriptor_write_waitrequest
	wire  [31:0] eth1_rx_dma_descriptor_write_address;                            // eth1_rx_dma:descriptor_write_address -> mm_interconnect_2:eth1_rx_dma_descriptor_write_address
	wire         eth1_rx_dma_descriptor_write_write;                              // eth1_rx_dma:descriptor_write_write -> mm_interconnect_2:eth1_rx_dma_descriptor_write_write
	wire  [31:0] eth1_rx_dma_descriptor_write_writedata;                          // eth1_rx_dma:descriptor_write_writedata -> mm_interconnect_2:eth1_rx_dma_descriptor_write_writedata
	wire         eth1_tx_dma_descriptor_write_waitrequest;                        // mm_interconnect_2:eth1_tx_dma_descriptor_write_waitrequest -> eth1_tx_dma:descriptor_write_waitrequest
	wire  [31:0] eth1_tx_dma_descriptor_write_address;                            // eth1_tx_dma:descriptor_write_address -> mm_interconnect_2:eth1_tx_dma_descriptor_write_address
	wire         eth1_tx_dma_descriptor_write_write;                              // eth1_tx_dma:descriptor_write_write -> mm_interconnect_2:eth1_tx_dma_descriptor_write_write
	wire  [31:0] eth1_tx_dma_descriptor_write_writedata;                          // eth1_tx_dma:descriptor_write_writedata -> mm_interconnect_2:eth1_tx_dma_descriptor_write_writedata
	wire         nios2_dma_descriptor_write_waitrequest;                          // mm_interconnect_2:nios2_dma_descriptor_write_waitrequest -> nios2_dma:descriptor_write_waitrequest
	wire  [31:0] nios2_dma_descriptor_write_address;                              // nios2_dma:descriptor_write_address -> mm_interconnect_2:nios2_dma_descriptor_write_address
	wire         nios2_dma_descriptor_write_write;                                // nios2_dma:descriptor_write_write -> mm_interconnect_2:nios2_dma_descriptor_write_write
	wire  [31:0] nios2_dma_descriptor_write_writedata;                            // nios2_dma:descriptor_write_writedata -> mm_interconnect_2:nios2_dma_descriptor_write_writedata
	wire  [31:0] eth0_tx_dma_m_read_readdata;                                     // mm_interconnect_2:eth0_tx_dma_m_read_readdata -> eth0_tx_dma:m_read_readdata
	wire         eth0_tx_dma_m_read_waitrequest;                                  // mm_interconnect_2:eth0_tx_dma_m_read_waitrequest -> eth0_tx_dma:m_read_waitrequest
	wire  [31:0] eth0_tx_dma_m_read_address;                                      // eth0_tx_dma:m_read_address -> mm_interconnect_2:eth0_tx_dma_m_read_address
	wire         eth0_tx_dma_m_read_read;                                         // eth0_tx_dma:m_read_read -> mm_interconnect_2:eth0_tx_dma_m_read_read
	wire         eth0_tx_dma_m_read_readdatavalid;                                // mm_interconnect_2:eth0_tx_dma_m_read_readdatavalid -> eth0_tx_dma:m_read_readdatavalid
	wire  [31:0] eth1_tx_dma_m_read_readdata;                                     // mm_interconnect_2:eth1_tx_dma_m_read_readdata -> eth1_tx_dma:m_read_readdata
	wire         eth1_tx_dma_m_read_waitrequest;                                  // mm_interconnect_2:eth1_tx_dma_m_read_waitrequest -> eth1_tx_dma:m_read_waitrequest
	wire  [31:0] eth1_tx_dma_m_read_address;                                      // eth1_tx_dma:m_read_address -> mm_interconnect_2:eth1_tx_dma_m_read_address
	wire         eth1_tx_dma_m_read_read;                                         // eth1_tx_dma:m_read_read -> mm_interconnect_2:eth1_tx_dma_m_read_read
	wire         eth1_tx_dma_m_read_readdatavalid;                                // mm_interconnect_2:eth1_tx_dma_m_read_readdatavalid -> eth1_tx_dma:m_read_readdatavalid
	wire         eth0_rx_dma_m_write_waitrequest;                                 // mm_interconnect_2:eth0_rx_dma_m_write_waitrequest -> eth0_rx_dma:m_write_waitrequest
	wire  [31:0] eth0_rx_dma_m_write_address;                                     // eth0_rx_dma:m_write_address -> mm_interconnect_2:eth0_rx_dma_m_write_address
	wire         eth0_rx_dma_m_write_write;                                       // eth0_rx_dma:m_write_write -> mm_interconnect_2:eth0_rx_dma_m_write_write
	wire   [7:0] eth0_rx_dma_m_write_writedata;                                   // eth0_rx_dma:m_write_writedata -> mm_interconnect_2:eth0_rx_dma_m_write_writedata
	wire         eth1_rx_dma_m_write_waitrequest;                                 // mm_interconnect_2:eth1_rx_dma_m_write_waitrequest -> eth1_rx_dma:m_write_waitrequest
	wire  [31:0] eth1_rx_dma_m_write_address;                                     // eth1_rx_dma:m_write_address -> mm_interconnect_2:eth1_rx_dma_m_write_address
	wire         eth1_rx_dma_m_write_write;                                       // eth1_rx_dma:m_write_write -> mm_interconnect_2:eth1_rx_dma_m_write_write
	wire   [7:0] eth1_rx_dma_m_write_writedata;                                   // eth1_rx_dma:m_write_writedata -> mm_interconnect_2:eth1_rx_dma_m_write_writedata
	wire         mm_interconnect_2_nios2_onchip_mem_s2_chipselect;                // mm_interconnect_2:nios2_onchip_mem_s2_chipselect -> nios2_onchip_mem:chipselect2
	wire  [31:0] mm_interconnect_2_nios2_onchip_mem_s2_readdata;                  // nios2_onchip_mem:readdata2 -> mm_interconnect_2:nios2_onchip_mem_s2_readdata
	wire  [15:0] mm_interconnect_2_nios2_onchip_mem_s2_address;                   // mm_interconnect_2:nios2_onchip_mem_s2_address -> nios2_onchip_mem:address2
	wire   [3:0] mm_interconnect_2_nios2_onchip_mem_s2_byteenable;                // mm_interconnect_2:nios2_onchip_mem_s2_byteenable -> nios2_onchip_mem:byteenable2
	wire         mm_interconnect_2_nios2_onchip_mem_s2_write;                     // mm_interconnect_2:nios2_onchip_mem_s2_write -> nios2_onchip_mem:write2
	wire  [31:0] mm_interconnect_2_nios2_onchip_mem_s2_writedata;                 // mm_interconnect_2:nios2_onchip_mem_s2_writedata -> nios2_onchip_mem:writedata2
	wire         mm_interconnect_2_nios2_onchip_mem_s2_clken;                     // mm_interconnect_2:nios2_onchip_mem_s2_clken -> nios2_onchip_mem:clken2
	wire         irq_mapper_receiver0_irq;                                        // eth0_rx_dma:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                        // eth0_tx_dma:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                        // eth1_rx_dma:csr_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                        // eth1_tx_dma:csr_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                        // nios2_dma:csr_irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                        // nios2_jtag_uart:av_irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                        // nios2_timer:irq -> irq_mapper:receiver6_irq
	wire  [31:0] nios2_cpu_irq_irq;                                               // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         irq_mapper_001_receiver0_irq;                                    // usb_jtag_uart:av_irq -> irq_mapper_001:receiver0_irq
	wire  [31:0] usb_nios2_cpu_irq_irq;                                           // irq_mapper_001:sender_irq -> usb_nios2_cpu:irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [audio_mem:reset, audio_position:reset_n, audio_position_end:reset_n, eth0_mdio:reset, eth0_rx_dma:system_reset_n, eth0_rx_fifo:out_reset_n, eth0_tx_dma:system_reset_n, eth0_tx_fifo:in_reset_n, eth1_mdio:reset, eth1_rx_dma:system_reset_n, eth1_rx_fifo:out_reset_n, eth1_tx_dma:system_reset_n, eth1_tx_fifo:in_reset_n, io_hex:reset_n, io_keys:reset_n, io_led_green:reset_n, io_led_red:reset_n, io_switches:reset_n, io_vga_sync:reset_n, mm_interconnect_0:nios2_dma_reset_reset_bridge_in_reset_reset, mm_interconnect_2:eth0_rx_dma_reset_reset_bridge_in_reset_reset, nios2_dma:system_reset_n, nios2_jtag_uart:rst_n, nios2_onchip_mem:reset, nios2_pll:reset, nios2_sysid:reset_n, nios2_timer:reset_n, sdram:reset_n, sram_multiplexer:RESET, usb_keycode:reset2, vga_background_offset:reset_n, vga_sprite_0:reset, vga_sprite_1:reset, vga_sprite_2:reset, vga_sprite_3:reset, vga_sprite_4:reset, vga_sprite_5:reset, vga_sprite_6:reset, vga_sprite_7:reset, vga_sprite_params:RESET]
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                          // rst_controller_001:reset_req -> [nios2_cpu:reset_req, rst_translator:reset_req_in]
	wire         nios2_cpu_debug_reset_request_reset;                             // nios2_cpu:debug_reset_request -> rst_controller_001:reset_in1
	wire         rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> [irq_mapper_001:reset, mm_interconnect_1:usb_nios2_cpu_reset_reset_bridge_in_reset_reset, rst_translator_001:in_reset, usb_hpi_address:reset_n, usb_hpi_cs:reset_n, usb_hpi_data:reset_n, usb_hpi_r:reset_n, usb_hpi_reset:reset_n, usb_hpi_w:reset_n, usb_jtag_uart:rst_n, usb_keycode:reset, usb_nios2_cpu:reset_n, usb_nios2_onchip_mem:reset, usb_nios2_sysid:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                          // rst_controller_002:reset_req -> [rst_translator_001:reset_req_in, usb_nios2_cpu:reset_req]

	ECE385_audio_mem audio_mem (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (mm_interconnect_0_audio_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_audio_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_audio_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_audio_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_audio_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_audio_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_audio_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.address2    (audio_mem_s2_address),                      //     s2.address
		.chipselect2 (audio_mem_s2_chipselect),                   //       .chipselect
		.clken2      (audio_mem_s2_clken),                        //       .clken
		.write2      (audio_mem_s2_write),                        //       .write
		.readdata2   (audio_mem_s2_readdata),                     //       .readdata
		.writedata2  (audio_mem_s2_writedata),                    //       .writedata
		.byteenable2 (audio_mem_s2_byteenable),                   //       .byteenable
		.clk2        (audio_mem_clk2_clk),                        //   clk2.clk
		.reset2      (audio_mem_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                      // (terminated)
		.freeze      (1'b0),                                      // (terminated)
		.reset_req2  (1'b0)                                       // (terminated)
	);

	ECE385_audio_position audio_position (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_audio_position_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_audio_position_s1_readdata), //                    .readdata
		.in_port  (audio_position_export)                         // external_connection.export
	);

	ECE385_audio_position_end audio_position_end (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_audio_position_end_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_audio_position_end_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_audio_position_end_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_audio_position_end_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_audio_position_end_s1_readdata),   //                    .readdata
		.out_port   (audio_position_end_export)                           // external_connection.export
	);

	lantian_mdio #(
		.CLOCK_DIVIDER (8'b00010100)
	) eth0_mdio (
		.avalon_slave_address     (mm_interconnect_0_eth0_mdio_avalon_slave_address),     // avalon_slave.address
		.avalon_slave_read        (mm_interconnect_0_eth0_mdio_avalon_slave_read),        //             .read
		.avalon_slave_readdata    (mm_interconnect_0_eth0_mdio_avalon_slave_readdata),    //             .readdata
		.avalon_slave_waitrequest (mm_interconnect_0_eth0_mdio_avalon_slave_waitrequest), //             .waitrequest
		.avalon_slave_write       (mm_interconnect_0_eth0_mdio_avalon_slave_write),       //             .write
		.avalon_slave_writedata   (mm_interconnect_0_eth0_mdio_avalon_slave_writedata),   //             .writedata
		.clk                      (clk_clk),                                              //        clock.clk
		.reset                    (rst_controller_reset_out_reset),                       //        reset.reset
		.mdc                      (eth0_mdio_mdc),                                        //         mdio.mdc
		.mdio_in                  (eth0_mdio_mdio_in),                                    //             .mdio_in
		.mdio_out                 (eth0_mdio_mdio_out),                                   //             .mdio_out
		.mdio_oen                 (eth0_mdio_mdio_oen),                                   //             .mdio_oen
		.phy_addr                 (eth0_mdio_phy_addr)                                    //             .phy_addr
	);

	ECE385_eth0_rx_dma eth0_rx_dma (
		.clk                           (clk_clk),                                      //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),              //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_eth0_rx_dma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_eth0_rx_dma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_eth0_rx_dma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_eth0_rx_dma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_eth0_rx_dma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_eth0_rx_dma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (eth0_rx_dma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (eth0_rx_dma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (eth0_rx_dma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (eth0_rx_dma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (eth0_rx_dma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (eth0_rx_dma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (eth0_rx_dma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (eth0_rx_dma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (eth0_rx_dma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                     //          csr_irq.irq
		.in_startofpacket              (eth0_rx_fifo_out_startofpacket),               //               in.startofpacket
		.in_endofpacket                (eth0_rx_fifo_out_endofpacket),                 //                 .endofpacket
		.in_data                       (eth0_rx_fifo_out_data),                        //                 .data
		.in_valid                      (eth0_rx_fifo_out_valid),                       //                 .valid
		.in_ready                      (eth0_rx_fifo_out_ready),                       //                 .ready
		.in_error                      (eth0_rx_fifo_out_error),                       //                 .error
		.m_write_waitrequest           (eth0_rx_dma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (eth0_rx_dma_m_write_address),                  //                 .address
		.m_write_write                 (eth0_rx_dma_m_write_write),                    //                 .write
		.m_write_writedata             (eth0_rx_dma_m_write_writedata)                 //                 .writedata
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (1024),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (3),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) eth0_rx_fifo (
		.in_clk            (eth0_rx_fifo_in_clk_clk),              //        in_clk.clk
		.in_reset_n        (eth0_rx_fifo_in_clk_reset_reset_n),    //  in_clk_reset.reset_n
		.out_clk           (clk_clk),                              //       out_clk.clk
		.out_reset_n       (~rst_controller_reset_out_reset),      // out_clk_reset.reset_n
		.in_data           (eth0_rx_fifo_in_data),                 //            in.data
		.in_valid          (eth0_rx_fifo_in_valid),                //              .valid
		.in_ready          (eth0_rx_fifo_in_ready),                //              .ready
		.in_startofpacket  (eth0_rx_fifo_in_startofpacket),        //              .startofpacket
		.in_endofpacket    (eth0_rx_fifo_in_endofpacket),          //              .endofpacket
		.in_error          (eth0_rx_fifo_in_error),                //              .error
		.out_data          (eth0_rx_fifo_out_data),                //           out.data
		.out_valid         (eth0_rx_fifo_out_valid),               //              .valid
		.out_ready         (eth0_rx_fifo_out_ready),               //              .ready
		.out_startofpacket (eth0_rx_fifo_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (eth0_rx_fifo_out_endofpacket),         //              .endofpacket
		.out_error         (eth0_rx_fifo_out_error),               //              .error
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_empty          (1'b0),                                 //   (terminated)
		.out_empty         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	ECE385_eth0_tx_dma eth0_tx_dma (
		.clk                           (clk_clk),                                      //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),              //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_eth0_tx_dma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_eth0_tx_dma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_eth0_tx_dma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_eth0_tx_dma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_eth0_tx_dma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_eth0_tx_dma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (eth0_tx_dma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (eth0_tx_dma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (eth0_tx_dma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (eth0_tx_dma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (eth0_tx_dma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (eth0_tx_dma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (eth0_tx_dma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (eth0_tx_dma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (eth0_tx_dma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                     //          csr_irq.irq
		.m_read_readdata               (eth0_tx_dma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (eth0_tx_dma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (eth0_tx_dma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (eth0_tx_dma_m_read_address),                   //                 .address
		.m_read_read                   (eth0_tx_dma_m_read_read),                      //                 .read
		.out_data                      (eth0_tx_dma_out_data),                         //              out.data
		.out_valid                     (eth0_tx_dma_out_valid),                        //                 .valid
		.out_ready                     (eth0_tx_dma_out_ready),                        //                 .ready
		.out_endofpacket               (eth0_tx_dma_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (eth0_tx_dma_out_startofpacket),                //                 .startofpacket
		.out_empty                     (eth0_tx_dma_out_empty)                         //                 .empty
	);

	ECE385_eth0_tx_dma_buffer #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) eth0_tx_dma_buffer (
		.in_clk_0_clk        (eth0_tx_dma_buffer_in_clk_0_clk),        // in_clk_0.clk
		.in_rst_0_reset      (eth0_tx_dma_buffer_in_rst_0_reset),      // in_rst_0.reset
		.in_0_data           (eth0_tx_dma_buffer_in_0_data),           //     in_0.data
		.in_0_valid          (eth0_tx_dma_buffer_in_0_valid),          //         .valid
		.in_0_ready          (eth0_tx_dma_buffer_in_0_ready),          //         .ready
		.in_0_startofpacket  (eth0_tx_dma_buffer_in_0_startofpacket),  //         .startofpacket
		.in_0_endofpacket    (eth0_tx_dma_buffer_in_0_endofpacket),    //         .endofpacket
		.in_0_empty          (eth0_tx_dma_buffer_in_0_empty),          //         .empty
		.out_0_data          (eth0_tx_dma_buffer_out_0_data),          //    out_0.data
		.out_0_valid         (eth0_tx_dma_buffer_out_0_valid),         //         .valid
		.out_0_ready         (eth0_tx_dma_buffer_out_0_ready),         //         .ready
		.out_0_startofpacket (eth0_tx_dma_buffer_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (eth0_tx_dma_buffer_out_0_endofpacket)    //         .endofpacket
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (4),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (1024),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) eth0_tx_fifo (
		.in_clk            (clk_clk),                              //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),      //  in_clk_reset.reset_n
		.out_clk           (eth0_tx_fifo_out_clk_clk),             //       out_clk.clk
		.out_reset_n       (eth0_tx_fifo_out_clk_reset_reset_n),   // out_clk_reset.reset_n
		.in_data           (eth0_tx_dma_out_data),                 //            in.data
		.in_valid          (eth0_tx_dma_out_valid),                //              .valid
		.in_ready          (eth0_tx_dma_out_ready),                //              .ready
		.in_startofpacket  (eth0_tx_dma_out_startofpacket),        //              .startofpacket
		.in_endofpacket    (eth0_tx_dma_out_endofpacket),          //              .endofpacket
		.in_empty          (eth0_tx_dma_out_empty),                //              .empty
		.out_data          (eth0_tx_fifo_out_data),                //           out.data
		.out_valid         (eth0_tx_fifo_out_valid),               //              .valid
		.out_ready         (eth0_tx_fifo_out_ready),               //              .ready
		.out_startofpacket (eth0_tx_fifo_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (eth0_tx_fifo_out_endofpacket),         //              .endofpacket
		.out_empty         (eth0_tx_fifo_out_empty),               //              .empty
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_error          (1'b0),                                 //   (terminated)
		.out_error         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	lantian_mdio #(
		.CLOCK_DIVIDER (8'b00010100)
	) eth1_mdio (
		.avalon_slave_address     (mm_interconnect_0_eth1_mdio_avalon_slave_address),     // avalon_slave.address
		.avalon_slave_read        (mm_interconnect_0_eth1_mdio_avalon_slave_read),        //             .read
		.avalon_slave_readdata    (mm_interconnect_0_eth1_mdio_avalon_slave_readdata),    //             .readdata
		.avalon_slave_waitrequest (mm_interconnect_0_eth1_mdio_avalon_slave_waitrequest), //             .waitrequest
		.avalon_slave_write       (mm_interconnect_0_eth1_mdio_avalon_slave_write),       //             .write
		.avalon_slave_writedata   (mm_interconnect_0_eth1_mdio_avalon_slave_writedata),   //             .writedata
		.clk                      (clk_clk),                                              //        clock.clk
		.reset                    (rst_controller_reset_out_reset),                       //        reset.reset
		.mdc                      (eth1_mdio_mdc),                                        //         mdio.mdc
		.mdio_in                  (eth1_mdio_mdio_in),                                    //             .mdio_in
		.mdio_out                 (eth1_mdio_mdio_out),                                   //             .mdio_out
		.mdio_oen                 (eth1_mdio_mdio_oen),                                   //             .mdio_oen
		.phy_addr                 (eth1_mdio_phy_addr)                                    //             .phy_addr
	);

	ECE385_eth0_rx_dma eth1_rx_dma (
		.clk                           (clk_clk),                                      //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),              //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_eth1_rx_dma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_eth1_rx_dma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_eth1_rx_dma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_eth1_rx_dma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_eth1_rx_dma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_eth1_rx_dma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (eth1_rx_dma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (eth1_rx_dma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (eth1_rx_dma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (eth1_rx_dma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (eth1_rx_dma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (eth1_rx_dma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (eth1_rx_dma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (eth1_rx_dma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (eth1_rx_dma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver2_irq),                     //          csr_irq.irq
		.in_startofpacket              (eth1_rx_fifo_out_startofpacket),               //               in.startofpacket
		.in_endofpacket                (eth1_rx_fifo_out_endofpacket),                 //                 .endofpacket
		.in_data                       (eth1_rx_fifo_out_data),                        //                 .data
		.in_valid                      (eth1_rx_fifo_out_valid),                       //                 .valid
		.in_ready                      (eth1_rx_fifo_out_ready),                       //                 .ready
		.in_error                      (eth1_rx_fifo_out_error),                       //                 .error
		.m_write_waitrequest           (eth1_rx_dma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (eth1_rx_dma_m_write_address),                  //                 .address
		.m_write_write                 (eth1_rx_dma_m_write_write),                    //                 .write
		.m_write_writedata             (eth1_rx_dma_m_write_writedata)                 //                 .writedata
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (1024),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (3),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) eth1_rx_fifo (
		.in_clk            (eth1_rx_fifo_in_clk_clk),              //        in_clk.clk
		.in_reset_n        (eth1_rx_fifo_in_clk_reset_reset_n),    //  in_clk_reset.reset_n
		.out_clk           (clk_clk),                              //       out_clk.clk
		.out_reset_n       (~rst_controller_reset_out_reset),      // out_clk_reset.reset_n
		.in_data           (eth1_rx_fifo_in_data),                 //            in.data
		.in_valid          (eth1_rx_fifo_in_valid),                //              .valid
		.in_ready          (eth1_rx_fifo_in_ready),                //              .ready
		.in_startofpacket  (eth1_rx_fifo_in_startofpacket),        //              .startofpacket
		.in_endofpacket    (eth1_rx_fifo_in_endofpacket),          //              .endofpacket
		.in_error          (eth1_rx_fifo_in_error),                //              .error
		.out_data          (eth1_rx_fifo_out_data),                //           out.data
		.out_valid         (eth1_rx_fifo_out_valid),               //              .valid
		.out_ready         (eth1_rx_fifo_out_ready),               //              .ready
		.out_startofpacket (eth1_rx_fifo_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (eth1_rx_fifo_out_endofpacket),         //              .endofpacket
		.out_error         (eth1_rx_fifo_out_error),               //              .error
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_empty          (1'b0),                                 //   (terminated)
		.out_empty         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	ECE385_eth1_tx_dma eth1_tx_dma (
		.clk                           (clk_clk),                                      //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),              //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_eth1_tx_dma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_eth1_tx_dma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_eth1_tx_dma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_eth1_tx_dma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_eth1_tx_dma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_eth1_tx_dma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (eth1_tx_dma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (eth1_tx_dma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (eth1_tx_dma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (eth1_tx_dma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (eth1_tx_dma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (eth1_tx_dma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (eth1_tx_dma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (eth1_tx_dma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (eth1_tx_dma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver3_irq),                     //          csr_irq.irq
		.m_read_readdata               (eth1_tx_dma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (eth1_tx_dma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (eth1_tx_dma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (eth1_tx_dma_m_read_address),                   //                 .address
		.m_read_read                   (eth1_tx_dma_m_read_read),                      //                 .read
		.out_data                      (eth1_tx_dma_out_data),                         //              out.data
		.out_valid                     (eth1_tx_dma_out_valid),                        //                 .valid
		.out_ready                     (eth1_tx_dma_out_ready),                        //                 .ready
		.out_endofpacket               (eth1_tx_dma_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (eth1_tx_dma_out_startofpacket),                //                 .startofpacket
		.out_empty                     (eth1_tx_dma_out_empty)                         //                 .empty
	);

	ECE385_eth0_tx_dma_buffer #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) eth1_tx_dma_buffer (
		.in_clk_0_clk        (eth1_tx_dma_buffer_in_clk_0_clk),        // in_clk_0.clk
		.in_rst_0_reset      (eth1_tx_dma_buffer_in_rst_0_reset),      // in_rst_0.reset
		.in_0_data           (eth1_tx_dma_buffer_in_0_data),           //     in_0.data
		.in_0_valid          (eth1_tx_dma_buffer_in_0_valid),          //         .valid
		.in_0_ready          (eth1_tx_dma_buffer_in_0_ready),          //         .ready
		.in_0_startofpacket  (eth1_tx_dma_buffer_in_0_startofpacket),  //         .startofpacket
		.in_0_endofpacket    (eth1_tx_dma_buffer_in_0_endofpacket),    //         .endofpacket
		.in_0_empty          (eth1_tx_dma_buffer_in_0_empty),          //         .empty
		.out_0_data          (eth1_tx_dma_buffer_out_0_data),          //    out_0.data
		.out_0_valid         (eth1_tx_dma_buffer_out_0_valid),         //         .valid
		.out_0_ready         (eth1_tx_dma_buffer_out_0_ready),         //         .ready
		.out_0_startofpacket (eth1_tx_dma_buffer_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (eth1_tx_dma_buffer_out_0_endofpacket)    //         .endofpacket
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (4),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (1024),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) eth1_tx_fifo (
		.in_clk            (clk_clk),                              //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),      //  in_clk_reset.reset_n
		.out_clk           (eth1_tx_fifo_out_clk_clk),             //       out_clk.clk
		.out_reset_n       (eth1_tx_fifo_out_clk_reset_reset_n),   // out_clk_reset.reset_n
		.in_data           (eth1_tx_dma_out_data),                 //            in.data
		.in_valid          (eth1_tx_dma_out_valid),                //              .valid
		.in_ready          (eth1_tx_dma_out_ready),                //              .ready
		.in_startofpacket  (eth1_tx_dma_out_startofpacket),        //              .startofpacket
		.in_endofpacket    (eth1_tx_dma_out_endofpacket),          //              .endofpacket
		.in_empty          (eth1_tx_dma_out_empty),                //              .empty
		.out_data          (eth1_tx_fifo_out_data),                //           out.data
		.out_valid         (eth1_tx_fifo_out_valid),               //              .valid
		.out_ready         (eth1_tx_fifo_out_ready),               //              .ready
		.out_startofpacket (eth1_tx_fifo_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (eth1_tx_fifo_out_endofpacket),         //              .endofpacket
		.out_empty         (eth1_tx_fifo_out_empty),               //              .empty
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_error          (1'b0),                                 //   (terminated)
		.out_error         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	ECE385_io_hex io_hex (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_io_hex_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_hex_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_hex_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_hex_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_hex_s1_readdata),   //                    .readdata
		.out_port   (io_hex_export)                           // external_connection.export
	);

	ECE385_io_keys io_keys (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_io_keys_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_io_keys_s1_readdata), //                    .readdata
		.in_port  (io_keys_export)                         // external_connection.export
	);

	ECE385_io_led_green io_led_green (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_io_led_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_led_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_led_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_led_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_led_green_s1_readdata),   //                    .readdata
		.out_port   (io_led_green_export)                           // external_connection.export
	);

	ECE385_io_led_red io_led_red (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_io_led_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_io_led_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_io_led_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_io_led_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_io_led_red_s1_readdata),   //                    .readdata
		.out_port   (io_led_red_export)                           // external_connection.export
	);

	ECE385_io_switches io_switches (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_io_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_io_switches_s1_readdata), //                    .readdata
		.in_port  (io_switches_export)                         // external_connection.export
	);

	ECE385_io_vga_sync io_vga_sync (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_io_vga_sync_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_io_vga_sync_s1_readdata), //                    .readdata
		.in_port  (io_vga_sync_export)                         // external_connection.export
	);

	ECE385_nios2_cpu nios2_cpu (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	ECE385_nios2_dma nios2_dma (
		.clk                           (clk_clk),                                    //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),            //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_nios2_dma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_nios2_dma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_nios2_dma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_nios2_dma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_nios2_dma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_nios2_dma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (nios2_dma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (nios2_dma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (nios2_dma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (nios2_dma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (nios2_dma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (nios2_dma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (nios2_dma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (nios2_dma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (nios2_dma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver4_irq),                   //          csr_irq.irq
		.m_read_readdata               (nios2_dma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (nios2_dma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (nios2_dma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (nios2_dma_m_read_address),                   //                 .address
		.m_read_read                   (nios2_dma_m_read_read),                      //                 .read
		.m_write_waitrequest           (nios2_dma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (nios2_dma_m_write_address),                  //                 .address
		.m_write_write                 (nios2_dma_m_write_write),                    //                 .write
		.m_write_writedata             (nios2_dma_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (nios2_dma_m_write_byteenable)                //                 .byteenable
	);

	ECE385_nios2_jtag_uart nios2_jtag_uart (
		.clk            (clk_clk),                                                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                 //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver5_irq)                                         //               irq.irq
	);

	ECE385_nios2_onchip_mem nios2_onchip_mem (
		.address     (mm_interconnect_0_nios2_onchip_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_nios2_onchip_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_nios2_onchip_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_nios2_onchip_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_nios2_onchip_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_nios2_onchip_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_nios2_onchip_mem_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_2_nios2_onchip_mem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_nios2_onchip_mem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_nios2_onchip_mem_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_nios2_onchip_mem_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_nios2_onchip_mem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_nios2_onchip_mem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_nios2_onchip_mem_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                                          //   clk1.clk
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.freeze      (1'b0),                                             // (terminated)
		.reset_req   (1'b0)                                              // (terminated)
	);

	ECE385_nios2_pll nios2_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read               (mm_interconnect_0_nios2_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_nios2_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_nios2_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_nios2_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_nios2_pll_pll_slave_writedata), //                      .writedata
		.inclk0             (clk_clk),                                         //                inclk0.clk
		.c0                 (nios2_pll_ethernet_clk),                          //                    c0.clk
		.c1                 (nios2_pll_sdram_clk),                             //                    c1.clk
		.c2                 (nios2_pll_c2_clk),                                //                    c2.clk
		.c3                 (nios2_pll_vga_clk),                               //                    c3.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (4'b0000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	ECE385_nios2_sysid nios2_sysid (
		.clock    (clk_clk),                                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //         reset.reset_n
		.readdata (mm_interconnect_0_nios2_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_nios2_sysid_control_slave_address)   //              .address
	);

	ECE385_nios2_timer nios2_timer (
		.clk        (clk_clk),                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             // reset.reset_n
		.address    (mm_interconnect_0_nios2_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_nios2_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_nios2_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_nios2_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_nios2_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)                     //   irq.irq
	);

	ECE385_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	SRAM_Multiplexer sram_multiplexer (
		.CLK           (clk_clk),                                          //  clock.clk
		.RESET         (rst_controller_reset_out_reset),                   //  reset.reset
		.AVL_READ      (mm_interconnect_0_sram_multiplexer_avl_read),      //    avl.read
		.AVL_WRITE     (mm_interconnect_0_sram_multiplexer_avl_write),     //       .write
		.AVL_WRITEDATA (mm_interconnect_0_sram_multiplexer_avl_writedata), //       .writedata
		.AVL_READDATA  (mm_interconnect_0_sram_multiplexer_avl_readdata),  //       .readdata
		.AVL_ADDR      (mm_interconnect_0_sram_multiplexer_avl_address),   //       .address
		.SRAM_ADDR     (sram_sram_addr),                                   //   sram.sram_addr
		.SRAM_CE_N     (sram_sram_ce_n),                                   //       .sram_ce_n
		.SRAM_DQ       (sram_sram_dq),                                     //       .sram_dq
		.SRAM_LB_N     (sram_sram_lb_n),                                   //       .sram_lb_n
		.SRAM_OE_N     (sram_sram_oe_n),                                   //       .sram_oe_n
		.SRAM_UB_N     (sram_sram_ub_n),                                   //       .sram_ub_n
		.SRAM_WE_N     (sram_sram_we_n),                                   //       .sram_we_n
		.VGA_DrawX     (vga_vga_drawx),                                    //    vga.vga_drawx
		.VGA_DrawY     (vga_vga_drawy),                                    //       .vga_drawy
		.VGA_VAL       (vga_vga_val),                                      //       .vga_val
		.CLK2          (nios2_pll_c2_clk)                                  // clock2.clk
	);

	ECE385_usb_hpi_address usb_hpi_address (
		.clk        (usb_clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_usb_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_usb_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_usb_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_usb_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_usb_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	ECE385_usb_hpi_cs usb_hpi_cs (
		.clk        (usb_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_usb_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_usb_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_usb_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_usb_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_usb_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	ECE385_usb_hpi_data usb_hpi_data (
		.clk        (usb_clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_1_usb_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_usb_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_usb_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_usb_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_usb_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	ECE385_usb_hpi_cs usb_hpi_r (
		.clk        (usb_clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_1_usb_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_usb_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_usb_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_usb_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_usb_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	ECE385_usb_hpi_cs usb_hpi_reset (
		.clk        (usb_clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_usb_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_usb_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_usb_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_usb_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_usb_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	ECE385_usb_hpi_cs usb_hpi_w (
		.clk        (usb_clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_1_usb_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_usb_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_usb_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_usb_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_usb_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	ECE385_nios2_jtag_uart usb_jtag_uart (
		.clk            (usb_clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                   //               irq.irq
	);

	ECE385_usb_keycode usb_keycode (
		.clk         (usb_clk_clk),                                 //   clk1.clk
		.address     (mm_interconnect_1_usb_keycode_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_usb_keycode_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_usb_keycode_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_usb_keycode_s1_write),      //       .write
		.readdata    (mm_interconnect_1_usb_keycode_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_usb_keycode_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_usb_keycode_s1_byteenable), //       .byteenable
		.reset       (rst_controller_002_reset_out_reset),          // reset1.reset
		.address2    (mm_interconnect_0_usb_keycode_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_usb_keycode_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_usb_keycode_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_usb_keycode_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_usb_keycode_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_usb_keycode_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_usb_keycode_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                     //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),              // reset2.reset
		.reset_req   (1'b0),                                        // (terminated)
		.freeze      (1'b0),                                        // (terminated)
		.reset_req2  (1'b0)                                         // (terminated)
	);

	ECE385_usb_nios2_cpu usb_nios2_cpu (
		.clk                                 (usb_clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (usb_nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (usb_nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (usb_nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (usb_nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (usb_nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (usb_nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (usb_nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (usb_nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (usb_nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (usb_nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (usb_nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (usb_nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (usb_nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                            //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       (usb_nios2_cpu_custom_instruction_master_readra)               // custom_instruction_master.readra
	);

	ECE385_usb_nios2_onchip_mem usb_nios2_onchip_mem (
		.clk        (usb_clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_1_usb_nios2_onchip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_usb_nios2_onchip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_usb_nios2_onchip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_usb_nios2_onchip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_1_usb_nios2_onchip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_usb_nios2_onchip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_usb_nios2_onchip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),                   // reset1.reset
		.reset_req  (1'b0),                                                 // (terminated)
		.freeze     (1'b0)                                                  // (terminated)
	);

	ECE385_nios2_sysid usb_nios2_sysid (
		.clock    (usb_clk_clk),                                              //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                      //         reset.reset_n
		.readdata (mm_interconnect_1_usb_nios2_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_usb_nios2_sysid_control_slave_address)   //              .address
	);

	ECE385_audio_position_end vga_background_offset (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_0_vga_background_offset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_vga_background_offset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_vga_background_offset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_vga_background_offset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_vga_background_offset_s1_readdata),   //                    .readdata
		.out_port   (vga_background_offset_export)                           // external_connection.export
	);

	ECE385_vga_sprite_0 vga_sprite_0 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_0_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_0_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_0_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_0_s2_clken),                        //       .clken
		.write2      (vga_sprite_0_s2_write),                        //       .write
		.readdata2   (vga_sprite_0_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_0_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_0_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_0_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_0_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	ECE385_vga_sprite_1 vga_sprite_1 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_1_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_1_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_1_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_1_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_1_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_1_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_1_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_1_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_1_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_1_s2_clken),                        //       .clken
		.write2      (vga_sprite_1_s2_write),                        //       .write
		.readdata2   (vga_sprite_1_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_1_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_1_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_1_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_1_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	ECE385_vga_sprite_2 vga_sprite_2 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_2_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_2_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_2_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_2_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_2_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_2_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_2_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_2_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_2_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_2_s2_clken),                        //       .clken
		.write2      (vga_sprite_2_s2_write),                        //       .write
		.readdata2   (vga_sprite_2_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_2_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_2_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_2_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_2_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	ECE385_vga_sprite_3 vga_sprite_3 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_3_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_3_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_3_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_3_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_3_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_3_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_3_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_3_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_3_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_3_s2_clken),                        //       .clken
		.write2      (vga_sprite_3_s2_write),                        //       .write
		.readdata2   (vga_sprite_3_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_3_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_3_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_3_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_3_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	ECE385_vga_sprite_4 vga_sprite_4 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_4_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_4_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_4_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_4_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_4_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_4_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_4_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_4_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_4_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_4_s2_clken),                        //       .clken
		.write2      (vga_sprite_4_s2_write),                        //       .write
		.readdata2   (vga_sprite_4_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_4_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_4_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_4_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_4_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	ECE385_vga_sprite_5 vga_sprite_5 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_5_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_5_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_5_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_5_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_5_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_5_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_5_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_5_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_5_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_5_s2_clken),                        //       .clken
		.write2      (vga_sprite_5_s2_write),                        //       .write
		.readdata2   (vga_sprite_5_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_5_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_5_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_5_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_5_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	ECE385_vga_sprite_6 vga_sprite_6 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_6_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_6_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_6_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_6_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_6_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_6_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_6_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_6_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_6_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_6_s2_clken),                        //       .clken
		.write2      (vga_sprite_6_s2_write),                        //       .write
		.readdata2   (vga_sprite_6_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_6_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_6_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_6_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_6_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	ECE385_vga_sprite_7 vga_sprite_7 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_vga_sprite_7_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_vga_sprite_7_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_vga_sprite_7_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_vga_sprite_7_s1_write),      //       .write
		.readdata    (mm_interconnect_0_vga_sprite_7_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_vga_sprite_7_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_vga_sprite_7_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.address2    (vga_sprite_7_s2_address),                      //     s2.address
		.chipselect2 (vga_sprite_7_s2_chipselect),                   //       .chipselect
		.clken2      (vga_sprite_7_s2_clken),                        //       .clken
		.write2      (vga_sprite_7_s2_write),                        //       .write
		.readdata2   (vga_sprite_7_s2_readdata),                     //       .readdata
		.writedata2  (vga_sprite_7_s2_writedata),                    //       .writedata
		.byteenable2 (vga_sprite_7_s2_byteenable),                   //       .byteenable
		.clk2        (vga_sprite_7_clk2_clk),                        //   clk2.clk
		.reset2      (vga_sprite_7_reset2_reset),                    // reset2.reset
		.reset_req   (1'b0),                                         // (terminated)
		.freeze      (1'b0),                                         // (terminated)
		.reset_req2  (1'b0)                                          // (terminated)
	);

	avalon_mm_passthrough #(
		.ADDR_WIDTH (8)
	) vga_sprite_params (
		.CLK            (clk_clk),                                           //        clock.clk
		.RESET          (rst_controller_reset_out_reset),                    //        reset.reset
		.AVL_READ       (mm_interconnect_0_vga_sprite_params_avl_read),      //          avl.read
		.AVL_WRITE      (mm_interconnect_0_vga_sprite_params_avl_write),     //             .write
		.AVL_WRITEDATA  (mm_interconnect_0_vga_sprite_params_avl_writedata), //             .writedata
		.AVL_READDATA   (mm_interconnect_0_vga_sprite_params_avl_readdata),  //             .readdata
		.AVL_ADDR       (mm_interconnect_0_vga_sprite_params_avl_address),   //             .address
		.PASS_CLK       (),                                                  // clock_source.clk
		.PASS_RESET     (vga_sprite_params_reset_reset),                     // reset_source.reset
		.PASS_ADDR      (vga_sprite_params_pass_address),                    //         pass.address
		.PASS_READ      (vga_sprite_params_pass_read),                       //             .read
		.PASS_READDATA  (vga_sprite_params_pass_readdata),                   //             .readdata
		.PASS_WRITE     (vga_sprite_params_pass_write),                      //             .write
		.PASS_WRITEDATA (vga_sprite_params_pass_writedata)                   //             .writedata
	);

	ECE385_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                                         //                             clk_0_clk.clk
		.nios2_cpu_reset_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),                              // nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_dma_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                                  // nios2_dma_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                 (nios2_cpu_data_master_address),                                   //                 nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest             (nios2_cpu_data_master_waitrequest),                               //                                      .waitrequest
		.nios2_cpu_data_master_byteenable              (nios2_cpu_data_master_byteenable),                                //                                      .byteenable
		.nios2_cpu_data_master_read                    (nios2_cpu_data_master_read),                                      //                                      .read
		.nios2_cpu_data_master_readdata                (nios2_cpu_data_master_readdata),                                  //                                      .readdata
		.nios2_cpu_data_master_write                   (nios2_cpu_data_master_write),                                     //                                      .write
		.nios2_cpu_data_master_writedata               (nios2_cpu_data_master_writedata),                                 //                                      .writedata
		.nios2_cpu_data_master_debugaccess             (nios2_cpu_data_master_debugaccess),                               //                                      .debugaccess
		.nios2_cpu_instruction_master_address          (nios2_cpu_instruction_master_address),                            //          nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest      (nios2_cpu_instruction_master_waitrequest),                        //                                      .waitrequest
		.nios2_cpu_instruction_master_read             (nios2_cpu_instruction_master_read),                               //                                      .read
		.nios2_cpu_instruction_master_readdata         (nios2_cpu_instruction_master_readdata),                           //                                      .readdata
		.nios2_dma_m_read_address                      (nios2_dma_m_read_address),                                        //                      nios2_dma_m_read.address
		.nios2_dma_m_read_waitrequest                  (nios2_dma_m_read_waitrequest),                                    //                                      .waitrequest
		.nios2_dma_m_read_read                         (nios2_dma_m_read_read),                                           //                                      .read
		.nios2_dma_m_read_readdata                     (nios2_dma_m_read_readdata),                                       //                                      .readdata
		.nios2_dma_m_read_readdatavalid                (nios2_dma_m_read_readdatavalid),                                  //                                      .readdatavalid
		.nios2_dma_m_write_address                     (nios2_dma_m_write_address),                                       //                     nios2_dma_m_write.address
		.nios2_dma_m_write_waitrequest                 (nios2_dma_m_write_waitrequest),                                   //                                      .waitrequest
		.nios2_dma_m_write_byteenable                  (nios2_dma_m_write_byteenable),                                    //                                      .byteenable
		.nios2_dma_m_write_write                       (nios2_dma_m_write_write),                                         //                                      .write
		.nios2_dma_m_write_writedata                   (nios2_dma_m_write_writedata),                                     //                                      .writedata
		.audio_mem_s1_address                          (mm_interconnect_0_audio_mem_s1_address),                          //                          audio_mem_s1.address
		.audio_mem_s1_write                            (mm_interconnect_0_audio_mem_s1_write),                            //                                      .write
		.audio_mem_s1_readdata                         (mm_interconnect_0_audio_mem_s1_readdata),                         //                                      .readdata
		.audio_mem_s1_writedata                        (mm_interconnect_0_audio_mem_s1_writedata),                        //                                      .writedata
		.audio_mem_s1_byteenable                       (mm_interconnect_0_audio_mem_s1_byteenable),                       //                                      .byteenable
		.audio_mem_s1_chipselect                       (mm_interconnect_0_audio_mem_s1_chipselect),                       //                                      .chipselect
		.audio_mem_s1_clken                            (mm_interconnect_0_audio_mem_s1_clken),                            //                                      .clken
		.audio_position_s1_address                     (mm_interconnect_0_audio_position_s1_address),                     //                     audio_position_s1.address
		.audio_position_s1_readdata                    (mm_interconnect_0_audio_position_s1_readdata),                    //                                      .readdata
		.audio_position_end_s1_address                 (mm_interconnect_0_audio_position_end_s1_address),                 //                 audio_position_end_s1.address
		.audio_position_end_s1_write                   (mm_interconnect_0_audio_position_end_s1_write),                   //                                      .write
		.audio_position_end_s1_readdata                (mm_interconnect_0_audio_position_end_s1_readdata),                //                                      .readdata
		.audio_position_end_s1_writedata               (mm_interconnect_0_audio_position_end_s1_writedata),               //                                      .writedata
		.audio_position_end_s1_chipselect              (mm_interconnect_0_audio_position_end_s1_chipselect),              //                                      .chipselect
		.eth0_mdio_avalon_slave_address                (mm_interconnect_0_eth0_mdio_avalon_slave_address),                //                eth0_mdio_avalon_slave.address
		.eth0_mdio_avalon_slave_write                  (mm_interconnect_0_eth0_mdio_avalon_slave_write),                  //                                      .write
		.eth0_mdio_avalon_slave_read                   (mm_interconnect_0_eth0_mdio_avalon_slave_read),                   //                                      .read
		.eth0_mdio_avalon_slave_readdata               (mm_interconnect_0_eth0_mdio_avalon_slave_readdata),               //                                      .readdata
		.eth0_mdio_avalon_slave_writedata              (mm_interconnect_0_eth0_mdio_avalon_slave_writedata),              //                                      .writedata
		.eth0_mdio_avalon_slave_waitrequest            (mm_interconnect_0_eth0_mdio_avalon_slave_waitrequest),            //                                      .waitrequest
		.eth0_rx_dma_csr_address                       (mm_interconnect_0_eth0_rx_dma_csr_address),                       //                       eth0_rx_dma_csr.address
		.eth0_rx_dma_csr_write                         (mm_interconnect_0_eth0_rx_dma_csr_write),                         //                                      .write
		.eth0_rx_dma_csr_read                          (mm_interconnect_0_eth0_rx_dma_csr_read),                          //                                      .read
		.eth0_rx_dma_csr_readdata                      (mm_interconnect_0_eth0_rx_dma_csr_readdata),                      //                                      .readdata
		.eth0_rx_dma_csr_writedata                     (mm_interconnect_0_eth0_rx_dma_csr_writedata),                     //                                      .writedata
		.eth0_rx_dma_csr_chipselect                    (mm_interconnect_0_eth0_rx_dma_csr_chipselect),                    //                                      .chipselect
		.eth0_tx_dma_csr_address                       (mm_interconnect_0_eth0_tx_dma_csr_address),                       //                       eth0_tx_dma_csr.address
		.eth0_tx_dma_csr_write                         (mm_interconnect_0_eth0_tx_dma_csr_write),                         //                                      .write
		.eth0_tx_dma_csr_read                          (mm_interconnect_0_eth0_tx_dma_csr_read),                          //                                      .read
		.eth0_tx_dma_csr_readdata                      (mm_interconnect_0_eth0_tx_dma_csr_readdata),                      //                                      .readdata
		.eth0_tx_dma_csr_writedata                     (mm_interconnect_0_eth0_tx_dma_csr_writedata),                     //                                      .writedata
		.eth0_tx_dma_csr_chipselect                    (mm_interconnect_0_eth0_tx_dma_csr_chipselect),                    //                                      .chipselect
		.eth1_mdio_avalon_slave_address                (mm_interconnect_0_eth1_mdio_avalon_slave_address),                //                eth1_mdio_avalon_slave.address
		.eth1_mdio_avalon_slave_write                  (mm_interconnect_0_eth1_mdio_avalon_slave_write),                  //                                      .write
		.eth1_mdio_avalon_slave_read                   (mm_interconnect_0_eth1_mdio_avalon_slave_read),                   //                                      .read
		.eth1_mdio_avalon_slave_readdata               (mm_interconnect_0_eth1_mdio_avalon_slave_readdata),               //                                      .readdata
		.eth1_mdio_avalon_slave_writedata              (mm_interconnect_0_eth1_mdio_avalon_slave_writedata),              //                                      .writedata
		.eth1_mdio_avalon_slave_waitrequest            (mm_interconnect_0_eth1_mdio_avalon_slave_waitrequest),            //                                      .waitrequest
		.eth1_rx_dma_csr_address                       (mm_interconnect_0_eth1_rx_dma_csr_address),                       //                       eth1_rx_dma_csr.address
		.eth1_rx_dma_csr_write                         (mm_interconnect_0_eth1_rx_dma_csr_write),                         //                                      .write
		.eth1_rx_dma_csr_read                          (mm_interconnect_0_eth1_rx_dma_csr_read),                          //                                      .read
		.eth1_rx_dma_csr_readdata                      (mm_interconnect_0_eth1_rx_dma_csr_readdata),                      //                                      .readdata
		.eth1_rx_dma_csr_writedata                     (mm_interconnect_0_eth1_rx_dma_csr_writedata),                     //                                      .writedata
		.eth1_rx_dma_csr_chipselect                    (mm_interconnect_0_eth1_rx_dma_csr_chipselect),                    //                                      .chipselect
		.eth1_tx_dma_csr_address                       (mm_interconnect_0_eth1_tx_dma_csr_address),                       //                       eth1_tx_dma_csr.address
		.eth1_tx_dma_csr_write                         (mm_interconnect_0_eth1_tx_dma_csr_write),                         //                                      .write
		.eth1_tx_dma_csr_read                          (mm_interconnect_0_eth1_tx_dma_csr_read),                          //                                      .read
		.eth1_tx_dma_csr_readdata                      (mm_interconnect_0_eth1_tx_dma_csr_readdata),                      //                                      .readdata
		.eth1_tx_dma_csr_writedata                     (mm_interconnect_0_eth1_tx_dma_csr_writedata),                     //                                      .writedata
		.eth1_tx_dma_csr_chipselect                    (mm_interconnect_0_eth1_tx_dma_csr_chipselect),                    //                                      .chipselect
		.io_hex_s1_address                             (mm_interconnect_0_io_hex_s1_address),                             //                             io_hex_s1.address
		.io_hex_s1_write                               (mm_interconnect_0_io_hex_s1_write),                               //                                      .write
		.io_hex_s1_readdata                            (mm_interconnect_0_io_hex_s1_readdata),                            //                                      .readdata
		.io_hex_s1_writedata                           (mm_interconnect_0_io_hex_s1_writedata),                           //                                      .writedata
		.io_hex_s1_chipselect                          (mm_interconnect_0_io_hex_s1_chipselect),                          //                                      .chipselect
		.io_keys_s1_address                            (mm_interconnect_0_io_keys_s1_address),                            //                            io_keys_s1.address
		.io_keys_s1_readdata                           (mm_interconnect_0_io_keys_s1_readdata),                           //                                      .readdata
		.io_led_green_s1_address                       (mm_interconnect_0_io_led_green_s1_address),                       //                       io_led_green_s1.address
		.io_led_green_s1_write                         (mm_interconnect_0_io_led_green_s1_write),                         //                                      .write
		.io_led_green_s1_readdata                      (mm_interconnect_0_io_led_green_s1_readdata),                      //                                      .readdata
		.io_led_green_s1_writedata                     (mm_interconnect_0_io_led_green_s1_writedata),                     //                                      .writedata
		.io_led_green_s1_chipselect                    (mm_interconnect_0_io_led_green_s1_chipselect),                    //                                      .chipselect
		.io_led_red_s1_address                         (mm_interconnect_0_io_led_red_s1_address),                         //                         io_led_red_s1.address
		.io_led_red_s1_write                           (mm_interconnect_0_io_led_red_s1_write),                           //                                      .write
		.io_led_red_s1_readdata                        (mm_interconnect_0_io_led_red_s1_readdata),                        //                                      .readdata
		.io_led_red_s1_writedata                       (mm_interconnect_0_io_led_red_s1_writedata),                       //                                      .writedata
		.io_led_red_s1_chipselect                      (mm_interconnect_0_io_led_red_s1_chipselect),                      //                                      .chipselect
		.io_switches_s1_address                        (mm_interconnect_0_io_switches_s1_address),                        //                        io_switches_s1.address
		.io_switches_s1_readdata                       (mm_interconnect_0_io_switches_s1_readdata),                       //                                      .readdata
		.io_vga_sync_s1_address                        (mm_interconnect_0_io_vga_sync_s1_address),                        //                        io_vga_sync_s1.address
		.io_vga_sync_s1_readdata                       (mm_interconnect_0_io_vga_sync_s1_readdata),                       //                                      .readdata
		.nios2_cpu_debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),             //             nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),               //                                      .write
		.nios2_cpu_debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),                //                                      .read
		.nios2_cpu_debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),            //                                      .readdata
		.nios2_cpu_debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),           //                                      .writedata
		.nios2_cpu_debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),          //                                      .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),         //                                      .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),         //                                      .debugaccess
		.nios2_dma_csr_address                         (mm_interconnect_0_nios2_dma_csr_address),                         //                         nios2_dma_csr.address
		.nios2_dma_csr_write                           (mm_interconnect_0_nios2_dma_csr_write),                           //                                      .write
		.nios2_dma_csr_read                            (mm_interconnect_0_nios2_dma_csr_read),                            //                                      .read
		.nios2_dma_csr_readdata                        (mm_interconnect_0_nios2_dma_csr_readdata),                        //                                      .readdata
		.nios2_dma_csr_writedata                       (mm_interconnect_0_nios2_dma_csr_writedata),                       //                                      .writedata
		.nios2_dma_csr_chipselect                      (mm_interconnect_0_nios2_dma_csr_chipselect),                      //                                      .chipselect
		.nios2_jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_address),     //     nios2_jtag_uart_avalon_jtag_slave.address
		.nios2_jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.nios2_jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.nios2_jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.nios2_jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.nios2_jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.nios2_jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_nios2_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.nios2_onchip_mem_s1_address                   (mm_interconnect_0_nios2_onchip_mem_s1_address),                   //                   nios2_onchip_mem_s1.address
		.nios2_onchip_mem_s1_write                     (mm_interconnect_0_nios2_onchip_mem_s1_write),                     //                                      .write
		.nios2_onchip_mem_s1_readdata                  (mm_interconnect_0_nios2_onchip_mem_s1_readdata),                  //                                      .readdata
		.nios2_onchip_mem_s1_writedata                 (mm_interconnect_0_nios2_onchip_mem_s1_writedata),                 //                                      .writedata
		.nios2_onchip_mem_s1_byteenable                (mm_interconnect_0_nios2_onchip_mem_s1_byteenable),                //                                      .byteenable
		.nios2_onchip_mem_s1_chipselect                (mm_interconnect_0_nios2_onchip_mem_s1_chipselect),                //                                      .chipselect
		.nios2_onchip_mem_s1_clken                     (mm_interconnect_0_nios2_onchip_mem_s1_clken),                     //                                      .clken
		.nios2_pll_pll_slave_address                   (mm_interconnect_0_nios2_pll_pll_slave_address),                   //                   nios2_pll_pll_slave.address
		.nios2_pll_pll_slave_write                     (mm_interconnect_0_nios2_pll_pll_slave_write),                     //                                      .write
		.nios2_pll_pll_slave_read                      (mm_interconnect_0_nios2_pll_pll_slave_read),                      //                                      .read
		.nios2_pll_pll_slave_readdata                  (mm_interconnect_0_nios2_pll_pll_slave_readdata),                  //                                      .readdata
		.nios2_pll_pll_slave_writedata                 (mm_interconnect_0_nios2_pll_pll_slave_writedata),                 //                                      .writedata
		.nios2_sysid_control_slave_address             (mm_interconnect_0_nios2_sysid_control_slave_address),             //             nios2_sysid_control_slave.address
		.nios2_sysid_control_slave_readdata            (mm_interconnect_0_nios2_sysid_control_slave_readdata),            //                                      .readdata
		.nios2_timer_s1_address                        (mm_interconnect_0_nios2_timer_s1_address),                        //                        nios2_timer_s1.address
		.nios2_timer_s1_write                          (mm_interconnect_0_nios2_timer_s1_write),                          //                                      .write
		.nios2_timer_s1_readdata                       (mm_interconnect_0_nios2_timer_s1_readdata),                       //                                      .readdata
		.nios2_timer_s1_writedata                      (mm_interconnect_0_nios2_timer_s1_writedata),                      //                                      .writedata
		.nios2_timer_s1_chipselect                     (mm_interconnect_0_nios2_timer_s1_chipselect),                     //                                      .chipselect
		.sdram_s1_address                              (mm_interconnect_0_sdram_s1_address),                              //                              sdram_s1.address
		.sdram_s1_write                                (mm_interconnect_0_sdram_s1_write),                                //                                      .write
		.sdram_s1_read                                 (mm_interconnect_0_sdram_s1_read),                                 //                                      .read
		.sdram_s1_readdata                             (mm_interconnect_0_sdram_s1_readdata),                             //                                      .readdata
		.sdram_s1_writedata                            (mm_interconnect_0_sdram_s1_writedata),                            //                                      .writedata
		.sdram_s1_byteenable                           (mm_interconnect_0_sdram_s1_byteenable),                           //                                      .byteenable
		.sdram_s1_readdatavalid                        (mm_interconnect_0_sdram_s1_readdatavalid),                        //                                      .readdatavalid
		.sdram_s1_waitrequest                          (mm_interconnect_0_sdram_s1_waitrequest),                          //                                      .waitrequest
		.sdram_s1_chipselect                           (mm_interconnect_0_sdram_s1_chipselect),                           //                                      .chipselect
		.sram_multiplexer_avl_address                  (mm_interconnect_0_sram_multiplexer_avl_address),                  //                  sram_multiplexer_avl.address
		.sram_multiplexer_avl_write                    (mm_interconnect_0_sram_multiplexer_avl_write),                    //                                      .write
		.sram_multiplexer_avl_read                     (mm_interconnect_0_sram_multiplexer_avl_read),                     //                                      .read
		.sram_multiplexer_avl_readdata                 (mm_interconnect_0_sram_multiplexer_avl_readdata),                 //                                      .readdata
		.sram_multiplexer_avl_writedata                (mm_interconnect_0_sram_multiplexer_avl_writedata),                //                                      .writedata
		.usb_keycode_s2_address                        (mm_interconnect_0_usb_keycode_s2_address),                        //                        usb_keycode_s2.address
		.usb_keycode_s2_write                          (mm_interconnect_0_usb_keycode_s2_write),                          //                                      .write
		.usb_keycode_s2_readdata                       (mm_interconnect_0_usb_keycode_s2_readdata),                       //                                      .readdata
		.usb_keycode_s2_writedata                      (mm_interconnect_0_usb_keycode_s2_writedata),                      //                                      .writedata
		.usb_keycode_s2_byteenable                     (mm_interconnect_0_usb_keycode_s2_byteenable),                     //                                      .byteenable
		.usb_keycode_s2_chipselect                     (mm_interconnect_0_usb_keycode_s2_chipselect),                     //                                      .chipselect
		.usb_keycode_s2_clken                          (mm_interconnect_0_usb_keycode_s2_clken),                          //                                      .clken
		.vga_background_offset_s1_address              (mm_interconnect_0_vga_background_offset_s1_address),              //              vga_background_offset_s1.address
		.vga_background_offset_s1_write                (mm_interconnect_0_vga_background_offset_s1_write),                //                                      .write
		.vga_background_offset_s1_readdata             (mm_interconnect_0_vga_background_offset_s1_readdata),             //                                      .readdata
		.vga_background_offset_s1_writedata            (mm_interconnect_0_vga_background_offset_s1_writedata),            //                                      .writedata
		.vga_background_offset_s1_chipselect           (mm_interconnect_0_vga_background_offset_s1_chipselect),           //                                      .chipselect
		.vga_sprite_0_s1_address                       (mm_interconnect_0_vga_sprite_0_s1_address),                       //                       vga_sprite_0_s1.address
		.vga_sprite_0_s1_write                         (mm_interconnect_0_vga_sprite_0_s1_write),                         //                                      .write
		.vga_sprite_0_s1_readdata                      (mm_interconnect_0_vga_sprite_0_s1_readdata),                      //                                      .readdata
		.vga_sprite_0_s1_writedata                     (mm_interconnect_0_vga_sprite_0_s1_writedata),                     //                                      .writedata
		.vga_sprite_0_s1_byteenable                    (mm_interconnect_0_vga_sprite_0_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_0_s1_chipselect                    (mm_interconnect_0_vga_sprite_0_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_0_s1_clken                         (mm_interconnect_0_vga_sprite_0_s1_clken),                         //                                      .clken
		.vga_sprite_1_s1_address                       (mm_interconnect_0_vga_sprite_1_s1_address),                       //                       vga_sprite_1_s1.address
		.vga_sprite_1_s1_write                         (mm_interconnect_0_vga_sprite_1_s1_write),                         //                                      .write
		.vga_sprite_1_s1_readdata                      (mm_interconnect_0_vga_sprite_1_s1_readdata),                      //                                      .readdata
		.vga_sprite_1_s1_writedata                     (mm_interconnect_0_vga_sprite_1_s1_writedata),                     //                                      .writedata
		.vga_sprite_1_s1_byteenable                    (mm_interconnect_0_vga_sprite_1_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_1_s1_chipselect                    (mm_interconnect_0_vga_sprite_1_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_1_s1_clken                         (mm_interconnect_0_vga_sprite_1_s1_clken),                         //                                      .clken
		.vga_sprite_2_s1_address                       (mm_interconnect_0_vga_sprite_2_s1_address),                       //                       vga_sprite_2_s1.address
		.vga_sprite_2_s1_write                         (mm_interconnect_0_vga_sprite_2_s1_write),                         //                                      .write
		.vga_sprite_2_s1_readdata                      (mm_interconnect_0_vga_sprite_2_s1_readdata),                      //                                      .readdata
		.vga_sprite_2_s1_writedata                     (mm_interconnect_0_vga_sprite_2_s1_writedata),                     //                                      .writedata
		.vga_sprite_2_s1_byteenable                    (mm_interconnect_0_vga_sprite_2_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_2_s1_chipselect                    (mm_interconnect_0_vga_sprite_2_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_2_s1_clken                         (mm_interconnect_0_vga_sprite_2_s1_clken),                         //                                      .clken
		.vga_sprite_3_s1_address                       (mm_interconnect_0_vga_sprite_3_s1_address),                       //                       vga_sprite_3_s1.address
		.vga_sprite_3_s1_write                         (mm_interconnect_0_vga_sprite_3_s1_write),                         //                                      .write
		.vga_sprite_3_s1_readdata                      (mm_interconnect_0_vga_sprite_3_s1_readdata),                      //                                      .readdata
		.vga_sprite_3_s1_writedata                     (mm_interconnect_0_vga_sprite_3_s1_writedata),                     //                                      .writedata
		.vga_sprite_3_s1_byteenable                    (mm_interconnect_0_vga_sprite_3_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_3_s1_chipselect                    (mm_interconnect_0_vga_sprite_3_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_3_s1_clken                         (mm_interconnect_0_vga_sprite_3_s1_clken),                         //                                      .clken
		.vga_sprite_4_s1_address                       (mm_interconnect_0_vga_sprite_4_s1_address),                       //                       vga_sprite_4_s1.address
		.vga_sprite_4_s1_write                         (mm_interconnect_0_vga_sprite_4_s1_write),                         //                                      .write
		.vga_sprite_4_s1_readdata                      (mm_interconnect_0_vga_sprite_4_s1_readdata),                      //                                      .readdata
		.vga_sprite_4_s1_writedata                     (mm_interconnect_0_vga_sprite_4_s1_writedata),                     //                                      .writedata
		.vga_sprite_4_s1_byteenable                    (mm_interconnect_0_vga_sprite_4_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_4_s1_chipselect                    (mm_interconnect_0_vga_sprite_4_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_4_s1_clken                         (mm_interconnect_0_vga_sprite_4_s1_clken),                         //                                      .clken
		.vga_sprite_5_s1_address                       (mm_interconnect_0_vga_sprite_5_s1_address),                       //                       vga_sprite_5_s1.address
		.vga_sprite_5_s1_write                         (mm_interconnect_0_vga_sprite_5_s1_write),                         //                                      .write
		.vga_sprite_5_s1_readdata                      (mm_interconnect_0_vga_sprite_5_s1_readdata),                      //                                      .readdata
		.vga_sprite_5_s1_writedata                     (mm_interconnect_0_vga_sprite_5_s1_writedata),                     //                                      .writedata
		.vga_sprite_5_s1_byteenable                    (mm_interconnect_0_vga_sprite_5_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_5_s1_chipselect                    (mm_interconnect_0_vga_sprite_5_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_5_s1_clken                         (mm_interconnect_0_vga_sprite_5_s1_clken),                         //                                      .clken
		.vga_sprite_6_s1_address                       (mm_interconnect_0_vga_sprite_6_s1_address),                       //                       vga_sprite_6_s1.address
		.vga_sprite_6_s1_write                         (mm_interconnect_0_vga_sprite_6_s1_write),                         //                                      .write
		.vga_sprite_6_s1_readdata                      (mm_interconnect_0_vga_sprite_6_s1_readdata),                      //                                      .readdata
		.vga_sprite_6_s1_writedata                     (mm_interconnect_0_vga_sprite_6_s1_writedata),                     //                                      .writedata
		.vga_sprite_6_s1_byteenable                    (mm_interconnect_0_vga_sprite_6_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_6_s1_chipselect                    (mm_interconnect_0_vga_sprite_6_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_6_s1_clken                         (mm_interconnect_0_vga_sprite_6_s1_clken),                         //                                      .clken
		.vga_sprite_7_s1_address                       (mm_interconnect_0_vga_sprite_7_s1_address),                       //                       vga_sprite_7_s1.address
		.vga_sprite_7_s1_write                         (mm_interconnect_0_vga_sprite_7_s1_write),                         //                                      .write
		.vga_sprite_7_s1_readdata                      (mm_interconnect_0_vga_sprite_7_s1_readdata),                      //                                      .readdata
		.vga_sprite_7_s1_writedata                     (mm_interconnect_0_vga_sprite_7_s1_writedata),                     //                                      .writedata
		.vga_sprite_7_s1_byteenable                    (mm_interconnect_0_vga_sprite_7_s1_byteenable),                    //                                      .byteenable
		.vga_sprite_7_s1_chipselect                    (mm_interconnect_0_vga_sprite_7_s1_chipselect),                    //                                      .chipselect
		.vga_sprite_7_s1_clken                         (mm_interconnect_0_vga_sprite_7_s1_clken),                         //                                      .clken
		.vga_sprite_params_avl_address                 (mm_interconnect_0_vga_sprite_params_avl_address),                 //                 vga_sprite_params_avl.address
		.vga_sprite_params_avl_write                   (mm_interconnect_0_vga_sprite_params_avl_write),                   //                                      .write
		.vga_sprite_params_avl_read                    (mm_interconnect_0_vga_sprite_params_avl_read),                    //                                      .read
		.vga_sprite_params_avl_readdata                (mm_interconnect_0_vga_sprite_params_avl_readdata),                //                                      .readdata
		.vga_sprite_params_avl_writedata               (mm_interconnect_0_vga_sprite_params_avl_writedata)                //                                      .writedata
	);

	ECE385_mm_interconnect_1 mm_interconnect_1 (
		.usb_clk_clk_clk                                 (usb_clk_clk),                                                   //                               usb_clk_clk.clk
		.usb_nios2_cpu_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                            // usb_nios2_cpu_reset_reset_bridge_in_reset.reset
		.usb_nios2_cpu_data_master_address               (usb_nios2_cpu_data_master_address),                             //                 usb_nios2_cpu_data_master.address
		.usb_nios2_cpu_data_master_waitrequest           (usb_nios2_cpu_data_master_waitrequest),                         //                                          .waitrequest
		.usb_nios2_cpu_data_master_byteenable            (usb_nios2_cpu_data_master_byteenable),                          //                                          .byteenable
		.usb_nios2_cpu_data_master_read                  (usb_nios2_cpu_data_master_read),                                //                                          .read
		.usb_nios2_cpu_data_master_readdata              (usb_nios2_cpu_data_master_readdata),                            //                                          .readdata
		.usb_nios2_cpu_data_master_write                 (usb_nios2_cpu_data_master_write),                               //                                          .write
		.usb_nios2_cpu_data_master_writedata             (usb_nios2_cpu_data_master_writedata),                           //                                          .writedata
		.usb_nios2_cpu_data_master_debugaccess           (usb_nios2_cpu_data_master_debugaccess),                         //                                          .debugaccess
		.usb_nios2_cpu_instruction_master_address        (usb_nios2_cpu_instruction_master_address),                      //          usb_nios2_cpu_instruction_master.address
		.usb_nios2_cpu_instruction_master_waitrequest    (usb_nios2_cpu_instruction_master_waitrequest),                  //                                          .waitrequest
		.usb_nios2_cpu_instruction_master_read           (usb_nios2_cpu_instruction_master_read),                         //                                          .read
		.usb_nios2_cpu_instruction_master_readdata       (usb_nios2_cpu_instruction_master_readdata),                     //                                          .readdata
		.usb_hpi_address_s1_address                      (mm_interconnect_1_usb_hpi_address_s1_address),                  //                        usb_hpi_address_s1.address
		.usb_hpi_address_s1_write                        (mm_interconnect_1_usb_hpi_address_s1_write),                    //                                          .write
		.usb_hpi_address_s1_readdata                     (mm_interconnect_1_usb_hpi_address_s1_readdata),                 //                                          .readdata
		.usb_hpi_address_s1_writedata                    (mm_interconnect_1_usb_hpi_address_s1_writedata),                //                                          .writedata
		.usb_hpi_address_s1_chipselect                   (mm_interconnect_1_usb_hpi_address_s1_chipselect),               //                                          .chipselect
		.usb_hpi_cs_s1_address                           (mm_interconnect_1_usb_hpi_cs_s1_address),                       //                             usb_hpi_cs_s1.address
		.usb_hpi_cs_s1_write                             (mm_interconnect_1_usb_hpi_cs_s1_write),                         //                                          .write
		.usb_hpi_cs_s1_readdata                          (mm_interconnect_1_usb_hpi_cs_s1_readdata),                      //                                          .readdata
		.usb_hpi_cs_s1_writedata                         (mm_interconnect_1_usb_hpi_cs_s1_writedata),                     //                                          .writedata
		.usb_hpi_cs_s1_chipselect                        (mm_interconnect_1_usb_hpi_cs_s1_chipselect),                    //                                          .chipselect
		.usb_hpi_data_s1_address                         (mm_interconnect_1_usb_hpi_data_s1_address),                     //                           usb_hpi_data_s1.address
		.usb_hpi_data_s1_write                           (mm_interconnect_1_usb_hpi_data_s1_write),                       //                                          .write
		.usb_hpi_data_s1_readdata                        (mm_interconnect_1_usb_hpi_data_s1_readdata),                    //                                          .readdata
		.usb_hpi_data_s1_writedata                       (mm_interconnect_1_usb_hpi_data_s1_writedata),                   //                                          .writedata
		.usb_hpi_data_s1_chipselect                      (mm_interconnect_1_usb_hpi_data_s1_chipselect),                  //                                          .chipselect
		.usb_hpi_r_s1_address                            (mm_interconnect_1_usb_hpi_r_s1_address),                        //                              usb_hpi_r_s1.address
		.usb_hpi_r_s1_write                              (mm_interconnect_1_usb_hpi_r_s1_write),                          //                                          .write
		.usb_hpi_r_s1_readdata                           (mm_interconnect_1_usb_hpi_r_s1_readdata),                       //                                          .readdata
		.usb_hpi_r_s1_writedata                          (mm_interconnect_1_usb_hpi_r_s1_writedata),                      //                                          .writedata
		.usb_hpi_r_s1_chipselect                         (mm_interconnect_1_usb_hpi_r_s1_chipselect),                     //                                          .chipselect
		.usb_hpi_reset_s1_address                        (mm_interconnect_1_usb_hpi_reset_s1_address),                    //                          usb_hpi_reset_s1.address
		.usb_hpi_reset_s1_write                          (mm_interconnect_1_usb_hpi_reset_s1_write),                      //                                          .write
		.usb_hpi_reset_s1_readdata                       (mm_interconnect_1_usb_hpi_reset_s1_readdata),                   //                                          .readdata
		.usb_hpi_reset_s1_writedata                      (mm_interconnect_1_usb_hpi_reset_s1_writedata),                  //                                          .writedata
		.usb_hpi_reset_s1_chipselect                     (mm_interconnect_1_usb_hpi_reset_s1_chipselect),                 //                                          .chipselect
		.usb_hpi_w_s1_address                            (mm_interconnect_1_usb_hpi_w_s1_address),                        //                              usb_hpi_w_s1.address
		.usb_hpi_w_s1_write                              (mm_interconnect_1_usb_hpi_w_s1_write),                          //                                          .write
		.usb_hpi_w_s1_readdata                           (mm_interconnect_1_usb_hpi_w_s1_readdata),                       //                                          .readdata
		.usb_hpi_w_s1_writedata                          (mm_interconnect_1_usb_hpi_w_s1_writedata),                      //                                          .writedata
		.usb_hpi_w_s1_chipselect                         (mm_interconnect_1_usb_hpi_w_s1_chipselect),                     //                                          .chipselect
		.usb_jtag_uart_avalon_jtag_slave_address         (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_address),     //           usb_jtag_uart_avalon_jtag_slave.address
		.usb_jtag_uart_avalon_jtag_slave_write           (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_write),       //                                          .write
		.usb_jtag_uart_avalon_jtag_slave_read            (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_read),        //                                          .read
		.usb_jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_readdata),    //                                          .readdata
		.usb_jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_writedata),   //                                          .writedata
		.usb_jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.usb_jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_1_usb_jtag_uart_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.usb_keycode_s1_address                          (mm_interconnect_1_usb_keycode_s1_address),                      //                            usb_keycode_s1.address
		.usb_keycode_s1_write                            (mm_interconnect_1_usb_keycode_s1_write),                        //                                          .write
		.usb_keycode_s1_readdata                         (mm_interconnect_1_usb_keycode_s1_readdata),                     //                                          .readdata
		.usb_keycode_s1_writedata                        (mm_interconnect_1_usb_keycode_s1_writedata),                    //                                          .writedata
		.usb_keycode_s1_byteenable                       (mm_interconnect_1_usb_keycode_s1_byteenable),                   //                                          .byteenable
		.usb_keycode_s1_chipselect                       (mm_interconnect_1_usb_keycode_s1_chipselect),                   //                                          .chipselect
		.usb_keycode_s1_clken                            (mm_interconnect_1_usb_keycode_s1_clken),                        //                                          .clken
		.usb_nios2_cpu_debug_mem_slave_address           (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_address),       //             usb_nios2_cpu_debug_mem_slave.address
		.usb_nios2_cpu_debug_mem_slave_write             (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_write),         //                                          .write
		.usb_nios2_cpu_debug_mem_slave_read              (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_read),          //                                          .read
		.usb_nios2_cpu_debug_mem_slave_readdata          (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_readdata),      //                                          .readdata
		.usb_nios2_cpu_debug_mem_slave_writedata         (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_writedata),     //                                          .writedata
		.usb_nios2_cpu_debug_mem_slave_byteenable        (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_byteenable),    //                                          .byteenable
		.usb_nios2_cpu_debug_mem_slave_waitrequest       (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_waitrequest),   //                                          .waitrequest
		.usb_nios2_cpu_debug_mem_slave_debugaccess       (mm_interconnect_1_usb_nios2_cpu_debug_mem_slave_debugaccess),   //                                          .debugaccess
		.usb_nios2_onchip_mem_s1_address                 (mm_interconnect_1_usb_nios2_onchip_mem_s1_address),             //                   usb_nios2_onchip_mem_s1.address
		.usb_nios2_onchip_mem_s1_write                   (mm_interconnect_1_usb_nios2_onchip_mem_s1_write),               //                                          .write
		.usb_nios2_onchip_mem_s1_readdata                (mm_interconnect_1_usb_nios2_onchip_mem_s1_readdata),            //                                          .readdata
		.usb_nios2_onchip_mem_s1_writedata               (mm_interconnect_1_usb_nios2_onchip_mem_s1_writedata),           //                                          .writedata
		.usb_nios2_onchip_mem_s1_byteenable              (mm_interconnect_1_usb_nios2_onchip_mem_s1_byteenable),          //                                          .byteenable
		.usb_nios2_onchip_mem_s1_chipselect              (mm_interconnect_1_usb_nios2_onchip_mem_s1_chipselect),          //                                          .chipselect
		.usb_nios2_onchip_mem_s1_clken                   (mm_interconnect_1_usb_nios2_onchip_mem_s1_clken),               //                                          .clken
		.usb_nios2_sysid_control_slave_address           (mm_interconnect_1_usb_nios2_sysid_control_slave_address),       //             usb_nios2_sysid_control_slave.address
		.usb_nios2_sysid_control_slave_readdata          (mm_interconnect_1_usb_nios2_sysid_control_slave_readdata)       //                                          .readdata
	);

	ECE385_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                 (clk_clk),                                          //                               clk_0_clk.clk
		.eth0_rx_dma_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // eth0_rx_dma_reset_reset_bridge_in_reset.reset
		.eth0_rx_dma_descriptor_read_address           (eth0_rx_dma_descriptor_read_address),              //             eth0_rx_dma_descriptor_read.address
		.eth0_rx_dma_descriptor_read_waitrequest       (eth0_rx_dma_descriptor_read_waitrequest),          //                                        .waitrequest
		.eth0_rx_dma_descriptor_read_read              (eth0_rx_dma_descriptor_read_read),                 //                                        .read
		.eth0_rx_dma_descriptor_read_readdata          (eth0_rx_dma_descriptor_read_readdata),             //                                        .readdata
		.eth0_rx_dma_descriptor_read_readdatavalid     (eth0_rx_dma_descriptor_read_readdatavalid),        //                                        .readdatavalid
		.eth0_rx_dma_descriptor_write_address          (eth0_rx_dma_descriptor_write_address),             //            eth0_rx_dma_descriptor_write.address
		.eth0_rx_dma_descriptor_write_waitrequest      (eth0_rx_dma_descriptor_write_waitrequest),         //                                        .waitrequest
		.eth0_rx_dma_descriptor_write_write            (eth0_rx_dma_descriptor_write_write),               //                                        .write
		.eth0_rx_dma_descriptor_write_writedata        (eth0_rx_dma_descriptor_write_writedata),           //                                        .writedata
		.eth0_rx_dma_m_write_address                   (eth0_rx_dma_m_write_address),                      //                     eth0_rx_dma_m_write.address
		.eth0_rx_dma_m_write_waitrequest               (eth0_rx_dma_m_write_waitrequest),                  //                                        .waitrequest
		.eth0_rx_dma_m_write_write                     (eth0_rx_dma_m_write_write),                        //                                        .write
		.eth0_rx_dma_m_write_writedata                 (eth0_rx_dma_m_write_writedata),                    //                                        .writedata
		.eth0_tx_dma_descriptor_read_address           (eth0_tx_dma_descriptor_read_address),              //             eth0_tx_dma_descriptor_read.address
		.eth0_tx_dma_descriptor_read_waitrequest       (eth0_tx_dma_descriptor_read_waitrequest),          //                                        .waitrequest
		.eth0_tx_dma_descriptor_read_read              (eth0_tx_dma_descriptor_read_read),                 //                                        .read
		.eth0_tx_dma_descriptor_read_readdata          (eth0_tx_dma_descriptor_read_readdata),             //                                        .readdata
		.eth0_tx_dma_descriptor_read_readdatavalid     (eth0_tx_dma_descriptor_read_readdatavalid),        //                                        .readdatavalid
		.eth0_tx_dma_descriptor_write_address          (eth0_tx_dma_descriptor_write_address),             //            eth0_tx_dma_descriptor_write.address
		.eth0_tx_dma_descriptor_write_waitrequest      (eth0_tx_dma_descriptor_write_waitrequest),         //                                        .waitrequest
		.eth0_tx_dma_descriptor_write_write            (eth0_tx_dma_descriptor_write_write),               //                                        .write
		.eth0_tx_dma_descriptor_write_writedata        (eth0_tx_dma_descriptor_write_writedata),           //                                        .writedata
		.eth0_tx_dma_m_read_address                    (eth0_tx_dma_m_read_address),                       //                      eth0_tx_dma_m_read.address
		.eth0_tx_dma_m_read_waitrequest                (eth0_tx_dma_m_read_waitrequest),                   //                                        .waitrequest
		.eth0_tx_dma_m_read_read                       (eth0_tx_dma_m_read_read),                          //                                        .read
		.eth0_tx_dma_m_read_readdata                   (eth0_tx_dma_m_read_readdata),                      //                                        .readdata
		.eth0_tx_dma_m_read_readdatavalid              (eth0_tx_dma_m_read_readdatavalid),                 //                                        .readdatavalid
		.eth1_rx_dma_descriptor_read_address           (eth1_rx_dma_descriptor_read_address),              //             eth1_rx_dma_descriptor_read.address
		.eth1_rx_dma_descriptor_read_waitrequest       (eth1_rx_dma_descriptor_read_waitrequest),          //                                        .waitrequest
		.eth1_rx_dma_descriptor_read_read              (eth1_rx_dma_descriptor_read_read),                 //                                        .read
		.eth1_rx_dma_descriptor_read_readdata          (eth1_rx_dma_descriptor_read_readdata),             //                                        .readdata
		.eth1_rx_dma_descriptor_read_readdatavalid     (eth1_rx_dma_descriptor_read_readdatavalid),        //                                        .readdatavalid
		.eth1_rx_dma_descriptor_write_address          (eth1_rx_dma_descriptor_write_address),             //            eth1_rx_dma_descriptor_write.address
		.eth1_rx_dma_descriptor_write_waitrequest      (eth1_rx_dma_descriptor_write_waitrequest),         //                                        .waitrequest
		.eth1_rx_dma_descriptor_write_write            (eth1_rx_dma_descriptor_write_write),               //                                        .write
		.eth1_rx_dma_descriptor_write_writedata        (eth1_rx_dma_descriptor_write_writedata),           //                                        .writedata
		.eth1_rx_dma_m_write_address                   (eth1_rx_dma_m_write_address),                      //                     eth1_rx_dma_m_write.address
		.eth1_rx_dma_m_write_waitrequest               (eth1_rx_dma_m_write_waitrequest),                  //                                        .waitrequest
		.eth1_rx_dma_m_write_write                     (eth1_rx_dma_m_write_write),                        //                                        .write
		.eth1_rx_dma_m_write_writedata                 (eth1_rx_dma_m_write_writedata),                    //                                        .writedata
		.eth1_tx_dma_descriptor_read_address           (eth1_tx_dma_descriptor_read_address),              //             eth1_tx_dma_descriptor_read.address
		.eth1_tx_dma_descriptor_read_waitrequest       (eth1_tx_dma_descriptor_read_waitrequest),          //                                        .waitrequest
		.eth1_tx_dma_descriptor_read_read              (eth1_tx_dma_descriptor_read_read),                 //                                        .read
		.eth1_tx_dma_descriptor_read_readdata          (eth1_tx_dma_descriptor_read_readdata),             //                                        .readdata
		.eth1_tx_dma_descriptor_read_readdatavalid     (eth1_tx_dma_descriptor_read_readdatavalid),        //                                        .readdatavalid
		.eth1_tx_dma_descriptor_write_address          (eth1_tx_dma_descriptor_write_address),             //            eth1_tx_dma_descriptor_write.address
		.eth1_tx_dma_descriptor_write_waitrequest      (eth1_tx_dma_descriptor_write_waitrequest),         //                                        .waitrequest
		.eth1_tx_dma_descriptor_write_write            (eth1_tx_dma_descriptor_write_write),               //                                        .write
		.eth1_tx_dma_descriptor_write_writedata        (eth1_tx_dma_descriptor_write_writedata),           //                                        .writedata
		.eth1_tx_dma_m_read_address                    (eth1_tx_dma_m_read_address),                       //                      eth1_tx_dma_m_read.address
		.eth1_tx_dma_m_read_waitrequest                (eth1_tx_dma_m_read_waitrequest),                   //                                        .waitrequest
		.eth1_tx_dma_m_read_read                       (eth1_tx_dma_m_read_read),                          //                                        .read
		.eth1_tx_dma_m_read_readdata                   (eth1_tx_dma_m_read_readdata),                      //                                        .readdata
		.eth1_tx_dma_m_read_readdatavalid              (eth1_tx_dma_m_read_readdatavalid),                 //                                        .readdatavalid
		.nios2_dma_descriptor_read_address             (nios2_dma_descriptor_read_address),                //               nios2_dma_descriptor_read.address
		.nios2_dma_descriptor_read_waitrequest         (nios2_dma_descriptor_read_waitrequest),            //                                        .waitrequest
		.nios2_dma_descriptor_read_read                (nios2_dma_descriptor_read_read),                   //                                        .read
		.nios2_dma_descriptor_read_readdata            (nios2_dma_descriptor_read_readdata),               //                                        .readdata
		.nios2_dma_descriptor_read_readdatavalid       (nios2_dma_descriptor_read_readdatavalid),          //                                        .readdatavalid
		.nios2_dma_descriptor_write_address            (nios2_dma_descriptor_write_address),               //              nios2_dma_descriptor_write.address
		.nios2_dma_descriptor_write_waitrequest        (nios2_dma_descriptor_write_waitrequest),           //                                        .waitrequest
		.nios2_dma_descriptor_write_write              (nios2_dma_descriptor_write_write),                 //                                        .write
		.nios2_dma_descriptor_write_writedata          (nios2_dma_descriptor_write_writedata),             //                                        .writedata
		.nios2_onchip_mem_s2_address                   (mm_interconnect_2_nios2_onchip_mem_s2_address),    //                     nios2_onchip_mem_s2.address
		.nios2_onchip_mem_s2_write                     (mm_interconnect_2_nios2_onchip_mem_s2_write),      //                                        .write
		.nios2_onchip_mem_s2_readdata                  (mm_interconnect_2_nios2_onchip_mem_s2_readdata),   //                                        .readdata
		.nios2_onchip_mem_s2_writedata                 (mm_interconnect_2_nios2_onchip_mem_s2_writedata),  //                                        .writedata
		.nios2_onchip_mem_s2_byteenable                (mm_interconnect_2_nios2_onchip_mem_s2_byteenable), //                                        .byteenable
		.nios2_onchip_mem_s2_chipselect                (mm_interconnect_2_nios2_onchip_mem_s2_chipselect), //                                        .chipselect
		.nios2_onchip_mem_s2_clken                     (mm_interconnect_2_nios2_onchip_mem_s2_clken)       //                                        .clken
	);

	ECE385_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.sender_irq    (nios2_cpu_irq_irq)                   //    sender.irq
	);

	ECE385_irq_mapper_001 irq_mapper_001 (
		.clk           (usb_clk_clk),                        //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.sender_irq    (usb_nios2_cpu_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~usb_reset_reset_n),                     // reset_in0.reset
		.clk            (usb_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
